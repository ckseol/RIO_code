function Bit#(300) encode(Bit#(300) x, Bit#(64) u);
	Bit#(300) y;
	y[0] = x[236]^x[238]^x[239]^x[241]^x[245]^x[255]^x[260]^x[264]^x[269]^x[271]^x[276]^x[279]^x[280]^x[285]^x[287]^x[289]^x[292]^x[293]^x[294]^x[295]^x[298]^u[63]^u[61]^u[60]^u[58]^u[54]^u[44]^u[39]^u[35]^u[30]^u[28]^u[23]^u[20]^u[19]^u[14]^u[12]^u[10]^u[7]^u[6]^u[5]^u[4]^u[1];
	y[1] = x[237]^x[239]^x[240]^x[242]^x[246]^x[256]^x[261]^x[265]^x[270]^x[272]^x[277]^x[280]^x[281]^x[286]^x[288]^x[290]^x[293]^x[294]^x[295]^x[296]^x[299]^u[62]^u[60]^u[59]^u[57]^u[53]^u[43]^u[38]^u[34]^u[29]^u[27]^u[22]^u[19]^u[18]^u[13]^u[11]^u[9]^u[6]^u[5]^u[4]^u[3]^u[0];
	y[2] = x[238]^x[240]^x[241]^x[243]^x[247]^x[257]^x[262]^x[266]^x[271]^x[273]^x[278]^x[281]^x[282]^x[287]^x[289]^x[291]^x[294]^x[295]^x[296]^x[297]^u[61]^u[59]^u[58]^u[56]^u[52]^u[42]^u[37]^u[33]^u[28]^u[26]^u[21]^u[18]^u[17]^u[12]^u[10]^u[8]^u[5]^u[4]^u[3]^u[2];
	y[3] = x[239]^x[241]^x[242]^x[244]^x[248]^x[258]^x[263]^x[267]^x[272]^x[274]^x[279]^x[282]^x[283]^x[288]^x[290]^x[292]^x[295]^x[296]^x[297]^x[298]^u[60]^u[58]^u[57]^u[55]^u[51]^u[41]^u[36]^u[32]^u[27]^u[25]^u[20]^u[17]^u[16]^u[11]^u[9]^u[7]^u[4]^u[3]^u[2]^u[1];
	y[4] = x[236]^x[238]^x[239]^x[240]^x[241]^x[242]^x[243]^x[249]^x[255]^x[259]^x[260]^x[268]^x[269]^x[271]^x[273]^x[275]^x[276]^x[279]^x[283]^x[284]^x[285]^x[287]^x[291]^x[292]^x[294]^x[295]^x[296]^x[297]^x[299]^u[63]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[50]^u[44]^u[40]^u[39]^u[31]^u[30]^u[28]^u[26]^u[24]^u[23]^u[20]^u[16]^u[15]^u[14]^u[12]^u[8]^u[7]^u[5]^u[4]^u[3]^u[2]^u[0];
	y[5] = x[237]^x[239]^x[240]^x[241]^x[242]^x[243]^x[244]^x[250]^x[256]^x[260]^x[261]^x[269]^x[270]^x[272]^x[274]^x[276]^x[277]^x[280]^x[284]^x[285]^x[286]^x[288]^x[292]^x[293]^x[295]^x[296]^x[297]^x[298]^u[62]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[49]^u[43]^u[39]^u[38]^u[30]^u[29]^u[27]^u[25]^u[23]^u[22]^u[19]^u[15]^u[14]^u[13]^u[11]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1];
	y[6] = x[236]^x[239]^x[240]^x[242]^x[243]^x[244]^x[251]^x[255]^x[257]^x[260]^x[261]^x[262]^x[264]^x[269]^x[270]^x[273]^x[275]^x[276]^x[277]^x[278]^x[279]^x[280]^x[281]^x[286]^x[292]^x[295]^x[296]^x[297]^x[299]^u[63]^u[60]^u[59]^u[57]^u[56]^u[55]^u[48]^u[44]^u[42]^u[39]^u[38]^u[37]^u[35]^u[30]^u[29]^u[26]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[13]^u[7]^u[4]^u[3]^u[2]^u[0];
	y[7] = x[237]^x[240]^x[241]^x[243]^x[244]^x[245]^x[252]^x[256]^x[258]^x[261]^x[262]^x[263]^x[265]^x[270]^x[271]^x[274]^x[276]^x[277]^x[278]^x[279]^x[280]^x[281]^x[282]^x[287]^x[293]^x[296]^x[297]^x[298]^u[62]^u[59]^u[58]^u[56]^u[55]^u[54]^u[47]^u[43]^u[41]^u[38]^u[37]^u[36]^u[34]^u[29]^u[28]^u[25]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[12]^u[6]^u[3]^u[2]^u[1];
	y[8] = x[236]^x[239]^x[242]^x[244]^x[246]^x[253]^x[255]^x[257]^x[259]^x[260]^x[262]^x[263]^x[266]^x[269]^x[272]^x[275]^x[276]^x[277]^x[278]^x[281]^x[282]^x[283]^x[285]^x[287]^x[288]^x[289]^x[292]^x[293]^x[295]^x[297]^x[299]^u[63]^u[60]^u[57]^u[55]^u[53]^u[46]^u[44]^u[42]^u[40]^u[39]^u[37]^u[36]^u[33]^u[30]^u[27]^u[24]^u[23]^u[22]^u[21]^u[18]^u[17]^u[16]^u[14]^u[12]^u[11]^u[10]^u[7]^u[6]^u[4]^u[2]^u[0];
	y[9] = x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[243]^x[247]^x[254]^x[255]^x[256]^x[258]^x[261]^x[263]^x[267]^x[269]^x[270]^x[271]^x[273]^x[277]^x[278]^x[280]^x[282]^x[283]^x[284]^x[285]^x[286]^x[287]^x[288]^x[290]^x[292]^x[295]^x[296]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[56]^u[52]^u[45]^u[44]^u[43]^u[41]^u[38]^u[36]^u[32]^u[30]^u[29]^u[28]^u[26]^u[22]^u[21]^u[19]^u[17]^u[16]^u[15]^u[14]^u[13]^u[12]^u[11]^u[9]^u[7]^u[4]^u[3];
	y[10] = x[236]^x[237]^x[240]^x[242]^x[244]^x[245]^x[248]^x[256]^x[257]^x[259]^x[260]^x[262]^x[268]^x[269]^x[270]^x[272]^x[274]^x[276]^x[278]^x[280]^x[281]^x[283]^x[284]^x[286]^x[288]^x[291]^x[292]^x[294]^x[295]^x[296]^x[297]^x[298]^u[63]^u[62]^u[59]^u[57]^u[55]^u[54]^u[51]^u[43]^u[42]^u[40]^u[39]^u[37]^u[31]^u[30]^u[29]^u[27]^u[25]^u[23]^u[21]^u[19]^u[18]^u[16]^u[15]^u[13]^u[11]^u[8]^u[7]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[11] = x[237]^x[238]^x[241]^x[243]^x[245]^x[246]^x[249]^x[257]^x[258]^x[260]^x[261]^x[263]^x[269]^x[270]^x[271]^x[273]^x[275]^x[277]^x[279]^x[281]^x[282]^x[284]^x[285]^x[287]^x[289]^x[292]^x[293]^x[295]^x[296]^x[297]^x[298]^x[299]^u[62]^u[61]^u[58]^u[56]^u[54]^u[53]^u[50]^u[42]^u[41]^u[39]^u[38]^u[36]^u[30]^u[29]^u[28]^u[26]^u[24]^u[22]^u[20]^u[18]^u[17]^u[15]^u[14]^u[12]^u[10]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[12] = x[238]^x[239]^x[242]^x[244]^x[246]^x[247]^x[250]^x[258]^x[259]^x[261]^x[262]^x[264]^x[270]^x[271]^x[272]^x[274]^x[276]^x[278]^x[280]^x[282]^x[283]^x[285]^x[286]^x[288]^x[290]^x[293]^x[294]^x[296]^x[297]^x[298]^x[299]^u[61]^u[60]^u[57]^u[55]^u[53]^u[52]^u[49]^u[41]^u[40]^u[38]^u[37]^u[35]^u[29]^u[28]^u[27]^u[25]^u[23]^u[21]^u[19]^u[17]^u[16]^u[14]^u[13]^u[11]^u[9]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[13] = x[236]^x[238]^x[240]^x[241]^x[243]^x[247]^x[248]^x[251]^x[255]^x[259]^x[262]^x[263]^x[264]^x[265]^x[269]^x[272]^x[273]^x[275]^x[276]^x[277]^x[280]^x[281]^x[283]^x[284]^x[285]^x[286]^x[291]^x[292]^x[293]^x[297]^x[299]^u[63]^u[61]^u[59]^u[58]^u[56]^u[52]^u[51]^u[48]^u[44]^u[40]^u[37]^u[36]^u[35]^u[34]^u[30]^u[27]^u[26]^u[24]^u[23]^u[22]^u[19]^u[18]^u[16]^u[15]^u[14]^u[13]^u[8]^u[7]^u[6]^u[2]^u[0];
	y[14] = x[236]^x[237]^x[238]^x[242]^x[244]^x[245]^x[248]^x[249]^x[252]^x[255]^x[256]^x[263]^x[265]^x[266]^x[269]^x[270]^x[271]^x[273]^x[274]^x[277]^x[278]^x[279]^x[280]^x[281]^x[282]^x[284]^x[286]^x[289]^x[295]^u[63]^u[62]^u[61]^u[57]^u[55]^u[54]^u[51]^u[50]^u[47]^u[44]^u[43]^u[36]^u[34]^u[33]^u[30]^u[29]^u[28]^u[26]^u[25]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[15]^u[13]^u[10]^u[4];
	y[15] = x[237]^x[238]^x[239]^x[243]^x[245]^x[246]^x[249]^x[250]^x[253]^x[256]^x[257]^x[264]^x[266]^x[267]^x[270]^x[271]^x[272]^x[274]^x[275]^x[278]^x[279]^x[280]^x[281]^x[282]^x[283]^x[285]^x[287]^x[290]^x[296]^u[62]^u[61]^u[60]^u[56]^u[54]^u[53]^u[50]^u[49]^u[46]^u[43]^u[42]^u[35]^u[33]^u[32]^u[29]^u[28]^u[27]^u[25]^u[24]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[14]^u[12]^u[9]^u[3];
	y[16] = x[238]^x[239]^x[240]^x[244]^x[246]^x[247]^x[250]^x[251]^x[254]^x[257]^x[258]^x[265]^x[267]^x[268]^x[271]^x[272]^x[273]^x[275]^x[276]^x[279]^x[280]^x[281]^x[282]^x[283]^x[284]^x[286]^x[288]^x[291]^x[297]^u[61]^u[60]^u[59]^u[55]^u[53]^u[52]^u[49]^u[48]^u[45]^u[42]^u[41]^u[34]^u[32]^u[31]^u[28]^u[27]^u[26]^u[24]^u[23]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[13]^u[11]^u[8]^u[2];
	y[17] = x[239]^x[240]^x[241]^x[245]^x[247]^x[248]^x[251]^x[252]^x[255]^x[258]^x[259]^x[266]^x[268]^x[269]^x[272]^x[273]^x[274]^x[276]^x[277]^x[280]^x[281]^x[282]^x[283]^x[284]^x[285]^x[287]^x[289]^x[292]^x[298]^u[60]^u[59]^u[58]^u[54]^u[52]^u[51]^u[48]^u[47]^u[44]^u[41]^u[40]^u[33]^u[31]^u[30]^u[27]^u[26]^u[25]^u[23]^u[22]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[10]^u[7]^u[1];
	y[18] = x[236]^x[238]^x[239]^x[240]^x[242]^x[245]^x[246]^x[248]^x[249]^x[252]^x[253]^x[255]^x[256]^x[259]^x[264]^x[267]^x[270]^x[271]^x[273]^x[274]^x[275]^x[276]^x[277]^x[278]^x[279]^x[280]^x[281]^x[282]^x[283]^x[284]^x[286]^x[287]^x[288]^x[289]^x[290]^x[292]^x[294]^x[295]^x[298]^x[299]^u[63]^u[61]^u[60]^u[59]^u[57]^u[54]^u[53]^u[51]^u[50]^u[47]^u[46]^u[44]^u[43]^u[40]^u[35]^u[32]^u[29]^u[28]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[9]^u[7]^u[5]^u[4]^u[1]^u[0];
	y[19] = x[237]^x[239]^x[240]^x[241]^x[243]^x[246]^x[247]^x[249]^x[250]^x[253]^x[254]^x[256]^x[257]^x[260]^x[265]^x[268]^x[271]^x[272]^x[274]^x[275]^x[276]^x[277]^x[278]^x[279]^x[280]^x[281]^x[282]^x[283]^x[284]^x[285]^x[287]^x[288]^x[289]^x[290]^x[291]^x[293]^x[295]^x[296]^x[299]^u[62]^u[60]^u[59]^u[58]^u[56]^u[53]^u[52]^u[50]^u[49]^u[46]^u[45]^u[43]^u[42]^u[39]^u[34]^u[31]^u[28]^u[27]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[8]^u[6]^u[4]^u[3]^u[0];
	y[20] = x[236]^x[239]^x[240]^x[242]^x[244]^x[245]^x[247]^x[248]^x[250]^x[251]^x[254]^x[257]^x[258]^x[260]^x[261]^x[264]^x[266]^x[271]^x[272]^x[273]^x[275]^x[277]^x[278]^x[281]^x[282]^x[283]^x[284]^x[286]^x[287]^x[288]^x[290]^x[291]^x[293]^x[295]^x[296]^x[297]^x[298]^u[63]^u[60]^u[59]^u[57]^u[55]^u[54]^u[52]^u[51]^u[49]^u[48]^u[45]^u[42]^u[41]^u[39]^u[38]^u[35]^u[33]^u[28]^u[27]^u[26]^u[24]^u[22]^u[21]^u[18]^u[17]^u[16]^u[15]^u[13]^u[12]^u[11]^u[9]^u[8]^u[6]^u[4]^u[3]^u[2]^u[1];
	y[21] = x[237]^x[240]^x[241]^x[243]^x[245]^x[246]^x[248]^x[249]^x[251]^x[252]^x[255]^x[258]^x[259]^x[261]^x[262]^x[265]^x[267]^x[272]^x[273]^x[274]^x[276]^x[278]^x[279]^x[282]^x[283]^x[284]^x[285]^x[287]^x[288]^x[289]^x[291]^x[292]^x[294]^x[296]^x[297]^x[298]^x[299]^u[62]^u[59]^u[58]^u[56]^u[54]^u[53]^u[51]^u[50]^u[48]^u[47]^u[44]^u[41]^u[40]^u[38]^u[37]^u[34]^u[32]^u[27]^u[26]^u[25]^u[23]^u[21]^u[20]^u[17]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[8]^u[7]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[22] = x[236]^x[239]^x[242]^x[244]^x[245]^x[246]^x[247]^x[249]^x[250]^x[252]^x[253]^x[255]^x[256]^x[259]^x[262]^x[263]^x[264]^x[266]^x[268]^x[269]^x[271]^x[273]^x[274]^x[275]^x[276]^x[277]^x[283]^x[284]^x[286]^x[287]^x[288]^x[290]^x[294]^x[297]^x[299]^u[63]^u[60]^u[57]^u[55]^u[54]^u[53]^u[52]^u[50]^u[49]^u[47]^u[46]^u[44]^u[43]^u[40]^u[37]^u[36]^u[35]^u[33]^u[31]^u[30]^u[28]^u[26]^u[25]^u[24]^u[23]^u[22]^u[16]^u[15]^u[13]^u[12]^u[11]^u[9]^u[5]^u[2]^u[0];
	y[23] = x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[243]^x[246]^x[247]^x[248]^x[250]^x[251]^x[253]^x[254]^x[255]^x[256]^x[257]^x[263]^x[265]^x[267]^x[270]^x[271]^x[272]^x[274]^x[275]^x[277]^x[278]^x[279]^x[280]^x[284]^x[288]^x[291]^x[292]^x[293]^x[294]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[56]^u[53]^u[52]^u[51]^u[49]^u[48]^u[46]^u[45]^u[44]^u[43]^u[42]^u[36]^u[34]^u[32]^u[29]^u[28]^u[27]^u[25]^u[24]^u[22]^u[21]^u[20]^u[19]^u[15]^u[11]^u[8]^u[7]^u[6]^u[5];
	y[24] = x[237]^x[238]^x[239]^x[240]^x[241]^x[242]^x[244]^x[247]^x[248]^x[249]^x[251]^x[252]^x[254]^x[255]^x[256]^x[257]^x[258]^x[264]^x[266]^x[268]^x[271]^x[272]^x[273]^x[275]^x[276]^x[278]^x[279]^x[280]^x[281]^x[285]^x[289]^x[292]^x[293]^x[294]^x[295]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[55]^u[52]^u[51]^u[50]^u[48]^u[47]^u[45]^u[44]^u[43]^u[42]^u[41]^u[35]^u[33]^u[31]^u[28]^u[27]^u[26]^u[24]^u[23]^u[21]^u[20]^u[19]^u[18]^u[14]^u[10]^u[7]^u[6]^u[5]^u[4];
	y[25] = x[236]^x[240]^x[242]^x[243]^x[248]^x[249]^x[250]^x[252]^x[253]^x[256]^x[257]^x[258]^x[259]^x[260]^x[264]^x[265]^x[267]^x[271]^x[272]^x[273]^x[274]^x[277]^x[281]^x[282]^x[285]^x[286]^x[287]^x[289]^x[290]^x[292]^x[296]^x[298]^u[63]^u[59]^u[57]^u[56]^u[51]^u[50]^u[49]^u[47]^u[46]^u[43]^u[42]^u[41]^u[40]^u[39]^u[35]^u[34]^u[32]^u[28]^u[27]^u[26]^u[25]^u[22]^u[18]^u[17]^u[14]^u[13]^u[12]^u[10]^u[9]^u[7]^u[3]^u[1];
	y[26] = x[236]^x[237]^x[238]^x[239]^x[243]^x[244]^x[245]^x[249]^x[250]^x[251]^x[253]^x[254]^x[255]^x[257]^x[258]^x[259]^x[261]^x[264]^x[265]^x[266]^x[268]^x[269]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[278]^x[279]^x[280]^x[282]^x[283]^x[285]^x[286]^x[288]^x[289]^x[290]^x[291]^x[292]^x[294]^x[295]^x[297]^x[298]^x[299]^u[63]^u[62]^u[61]^u[60]^u[56]^u[55]^u[54]^u[50]^u[49]^u[48]^u[46]^u[45]^u[44]^u[42]^u[41]^u[40]^u[38]^u[35]^u[34]^u[33]^u[31]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[21]^u[20]^u[19]^u[17]^u[16]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[27] = x[236]^x[237]^x[240]^x[241]^x[244]^x[246]^x[250]^x[251]^x[252]^x[254]^x[256]^x[258]^x[259]^x[262]^x[264]^x[265]^x[266]^x[267]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[277]^x[281]^x[283]^x[284]^x[285]^x[286]^x[290]^x[291]^x[294]^x[296]^x[299]^u[63]^u[62]^u[59]^u[58]^u[55]^u[53]^u[49]^u[48]^u[47]^u[45]^u[43]^u[41]^u[40]^u[37]^u[35]^u[34]^u[33]^u[32]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[22]^u[18]^u[16]^u[15]^u[14]^u[13]^u[9]^u[8]^u[5]^u[3]^u[0];
	y[28] = x[236]^x[237]^x[239]^x[242]^x[247]^x[251]^x[252]^x[253]^x[257]^x[259]^x[263]^x[264]^x[265]^x[266]^x[267]^x[268]^x[269]^x[272]^x[273]^x[274]^x[275]^x[278]^x[279]^x[280]^x[282]^x[284]^x[286]^x[289]^x[291]^x[293]^x[294]^x[297]^x[298]^u[63]^u[62]^u[60]^u[57]^u[52]^u[48]^u[47]^u[46]^u[42]^u[40]^u[36]^u[35]^u[34]^u[33]^u[32]^u[31]^u[30]^u[27]^u[26]^u[25]^u[24]^u[21]^u[20]^u[19]^u[17]^u[15]^u[13]^u[10]^u[8]^u[6]^u[5]^u[2]^u[1];
	y[29] = x[237]^x[238]^x[240]^x[243]^x[248]^x[252]^x[253]^x[254]^x[258]^x[260]^x[264]^x[265]^x[266]^x[267]^x[268]^x[269]^x[270]^x[273]^x[274]^x[275]^x[276]^x[279]^x[280]^x[281]^x[283]^x[285]^x[287]^x[290]^x[292]^x[294]^x[295]^x[298]^x[299]^u[62]^u[61]^u[59]^u[56]^u[51]^u[47]^u[46]^u[45]^u[41]^u[39]^u[35]^u[34]^u[33]^u[32]^u[31]^u[30]^u[29]^u[26]^u[25]^u[24]^u[23]^u[20]^u[19]^u[18]^u[16]^u[14]^u[12]^u[9]^u[7]^u[5]^u[4]^u[1]^u[0];
	y[30] = x[236]^x[244]^x[245]^x[249]^x[253]^x[254]^x[259]^x[260]^x[261]^x[264]^x[265]^x[266]^x[267]^x[268]^x[270]^x[274]^x[275]^x[277]^x[279]^x[281]^x[282]^x[284]^x[285]^x[286]^x[287]^x[288]^x[289]^x[291]^x[292]^x[294]^x[296]^x[298]^x[299]^u[63]^u[55]^u[54]^u[50]^u[46]^u[45]^u[40]^u[39]^u[38]^u[35]^u[34]^u[33]^u[32]^u[31]^u[29]^u[25]^u[24]^u[22]^u[20]^u[18]^u[17]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[8]^u[7]^u[5]^u[3]^u[1]^u[0];
	y[31] = x[236]^x[237]^x[238]^x[239]^x[241]^x[246]^x[250]^x[254]^x[261]^x[262]^x[264]^x[265]^x[266]^x[267]^x[268]^x[275]^x[278]^x[279]^x[282]^x[283]^x[286]^x[288]^x[290]^x[294]^x[297]^x[298]^x[299]^u[63]^u[62]^u[61]^u[60]^u[58]^u[53]^u[49]^u[45]^u[38]^u[37]^u[35]^u[34]^u[33]^u[32]^u[31]^u[24]^u[21]^u[20]^u[17]^u[16]^u[13]^u[11]^u[9]^u[5]^u[2]^u[1]^u[0];
	y[32] = x[236]^x[237]^x[240]^x[241]^x[242]^x[245]^x[247]^x[251]^x[260]^x[262]^x[263]^x[264]^x[265]^x[266]^x[267]^x[268]^x[271]^x[283]^x[284]^x[285]^x[291]^x[292]^x[293]^x[294]^x[299]^u[63]^u[62]^u[59]^u[58]^u[57]^u[54]^u[52]^u[48]^u[39]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32]^u[31]^u[28]^u[16]^u[15]^u[14]^u[8]^u[7]^u[6]^u[5]^u[0];
	y[33] = x[236]^x[237]^x[239]^x[242]^x[243]^x[245]^x[246]^x[248]^x[252]^x[255]^x[260]^x[261]^x[263]^x[265]^x[266]^x[267]^x[268]^x[271]^x[272]^x[276]^x[279]^x[280]^x[284]^x[286]^x[287]^x[289]^x[298]^u[63]^u[62]^u[60]^u[57]^u[56]^u[54]^u[53]^u[51]^u[47]^u[44]^u[39]^u[38]^u[36]^u[34]^u[33]^u[32]^u[31]^u[28]^u[27]^u[23]^u[20]^u[19]^u[15]^u[13]^u[12]^u[10]^u[1];
	y[34] = x[237]^x[238]^x[240]^x[243]^x[244]^x[246]^x[247]^x[249]^x[253]^x[256]^x[261]^x[262]^x[264]^x[266]^x[267]^x[268]^x[269]^x[272]^x[273]^x[277]^x[280]^x[281]^x[285]^x[287]^x[288]^x[290]^x[299]^u[62]^u[61]^u[59]^u[56]^u[55]^u[53]^u[52]^u[50]^u[46]^u[43]^u[38]^u[37]^u[35]^u[33]^u[32]^u[31]^u[30]^u[27]^u[26]^u[22]^u[19]^u[18]^u[14]^u[12]^u[11]^u[9]^u[0];
	y[35] = x[236]^x[244]^x[247]^x[248]^x[250]^x[254]^x[255]^x[257]^x[260]^x[262]^x[263]^x[264]^x[265]^x[267]^x[268]^x[270]^x[271]^x[273]^x[274]^x[276]^x[278]^x[279]^x[280]^x[281]^x[282]^x[285]^x[286]^x[287]^x[288]^x[291]^x[292]^x[293]^x[294]^x[295]^x[298]^u[63]^u[55]^u[52]^u[51]^u[49]^u[45]^u[44]^u[42]^u[39]^u[37]^u[36]^u[35]^u[34]^u[32]^u[31]^u[29]^u[28]^u[26]^u[25]^u[23]^u[21]^u[20]^u[19]^u[18]^u[17]^u[14]^u[13]^u[12]^u[11]^u[8]^u[7]^u[6]^u[5]^u[4]^u[1];
	y[36] = x[237]^x[245]^x[248]^x[249]^x[251]^x[255]^x[256]^x[258]^x[261]^x[263]^x[264]^x[265]^x[266]^x[268]^x[269]^x[271]^x[272]^x[274]^x[275]^x[277]^x[279]^x[280]^x[281]^x[282]^x[283]^x[286]^x[287]^x[288]^x[289]^x[292]^x[293]^x[294]^x[295]^x[296]^x[299]^u[62]^u[54]^u[51]^u[50]^u[48]^u[44]^u[43]^u[41]^u[38]^u[36]^u[35]^u[34]^u[33]^u[31]^u[30]^u[28]^u[27]^u[25]^u[24]^u[22]^u[20]^u[19]^u[18]^u[17]^u[16]^u[13]^u[12]^u[11]^u[10]^u[7]^u[6]^u[5]^u[4]^u[3]^u[0];
	y[37] = x[236]^x[239]^x[241]^x[245]^x[246]^x[249]^x[250]^x[252]^x[255]^x[256]^x[257]^x[259]^x[260]^x[262]^x[265]^x[266]^x[267]^x[270]^x[271]^x[272]^x[273]^x[275]^x[278]^x[279]^x[281]^x[282]^x[283]^x[284]^x[285]^x[288]^x[290]^x[292]^x[296]^x[297]^x[298]^u[63]^u[60]^u[58]^u[54]^u[53]^u[50]^u[49]^u[47]^u[44]^u[43]^u[42]^u[40]^u[39]^u[37]^u[34]^u[33]^u[32]^u[29]^u[28]^u[27]^u[26]^u[24]^u[21]^u[20]^u[18]^u[17]^u[16]^u[15]^u[14]^u[11]^u[9]^u[7]^u[3]^u[2]^u[1];
	y[38] = x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[242]^x[245]^x[246]^x[247]^x[250]^x[251]^x[253]^x[255]^x[256]^x[257]^x[258]^x[261]^x[263]^x[264]^x[266]^x[267]^x[268]^x[269]^x[272]^x[273]^x[274]^x[282]^x[283]^x[284]^x[286]^x[287]^x[291]^x[292]^x[294]^x[295]^x[297]^x[299]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[54]^u[53]^u[52]^u[49]^u[48]^u[46]^u[44]^u[43]^u[42]^u[41]^u[38]^u[36]^u[35]^u[33]^u[32]^u[31]^u[30]^u[27]^u[26]^u[25]^u[17]^u[16]^u[15]^u[13]^u[12]^u[8]^u[7]^u[5]^u[4]^u[2]^u[0];
	y[39] = x[237]^x[238]^x[239]^x[240]^x[241]^x[242]^x[243]^x[246]^x[247]^x[248]^x[251]^x[252]^x[254]^x[256]^x[257]^x[258]^x[259]^x[262]^x[264]^x[265]^x[267]^x[268]^x[269]^x[270]^x[273]^x[274]^x[275]^x[283]^x[284]^x[285]^x[287]^x[288]^x[292]^x[293]^x[295]^x[296]^x[298]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[53]^u[52]^u[51]^u[48]^u[47]^u[45]^u[43]^u[42]^u[41]^u[40]^u[37]^u[35]^u[34]^u[32]^u[31]^u[30]^u[29]^u[26]^u[25]^u[24]^u[16]^u[15]^u[14]^u[12]^u[11]^u[7]^u[6]^u[4]^u[3]^u[1];
	y[40] = x[238]^x[239]^x[240]^x[241]^x[242]^x[243]^x[244]^x[247]^x[248]^x[249]^x[252]^x[253]^x[255]^x[257]^x[258]^x[259]^x[260]^x[263]^x[265]^x[266]^x[268]^x[269]^x[270]^x[271]^x[274]^x[275]^x[276]^x[284]^x[285]^x[286]^x[288]^x[289]^x[293]^x[294]^x[296]^x[297]^x[299]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[52]^u[51]^u[50]^u[47]^u[46]^u[44]^u[42]^u[41]^u[40]^u[39]^u[36]^u[34]^u[33]^u[31]^u[30]^u[29]^u[28]^u[25]^u[24]^u[23]^u[15]^u[14]^u[13]^u[11]^u[10]^u[6]^u[5]^u[3]^u[2]^u[0];
	y[41] = x[236]^x[238]^x[240]^x[242]^x[243]^x[244]^x[248]^x[249]^x[250]^x[253]^x[254]^x[255]^x[256]^x[258]^x[259]^x[261]^x[266]^x[267]^x[270]^x[272]^x[275]^x[277]^x[279]^x[280]^x[286]^x[290]^x[292]^x[293]^x[297]^u[63]^u[61]^u[59]^u[57]^u[56]^u[55]^u[51]^u[50]^u[49]^u[46]^u[45]^u[44]^u[43]^u[41]^u[40]^u[38]^u[33]^u[32]^u[29]^u[27]^u[24]^u[22]^u[20]^u[19]^u[13]^u[9]^u[7]^u[6]^u[2];
	y[42] = x[237]^x[239]^x[241]^x[243]^x[244]^x[245]^x[249]^x[250]^x[251]^x[254]^x[255]^x[256]^x[257]^x[259]^x[260]^x[262]^x[267]^x[268]^x[271]^x[273]^x[276]^x[278]^x[280]^x[281]^x[287]^x[291]^x[293]^x[294]^x[298]^u[62]^u[60]^u[58]^u[56]^u[55]^u[54]^u[50]^u[49]^u[48]^u[45]^u[44]^u[43]^u[42]^u[40]^u[39]^u[37]^u[32]^u[31]^u[28]^u[26]^u[23]^u[21]^u[19]^u[18]^u[12]^u[8]^u[6]^u[5]^u[1];
	y[43] = x[236]^x[239]^x[240]^x[241]^x[242]^x[244]^x[246]^x[250]^x[251]^x[252]^x[256]^x[257]^x[258]^x[261]^x[263]^x[264]^x[268]^x[271]^x[272]^x[274]^x[276]^x[277]^x[280]^x[281]^x[282]^x[285]^x[287]^x[288]^x[289]^x[293]^x[298]^x[299]^u[63]^u[60]^u[59]^u[58]^u[57]^u[55]^u[53]^u[49]^u[48]^u[47]^u[43]^u[42]^u[41]^u[38]^u[36]^u[35]^u[31]^u[28]^u[27]^u[25]^u[23]^u[22]^u[19]^u[18]^u[17]^u[14]^u[12]^u[11]^u[10]^u[6]^u[1]^u[0];
	y[44] = x[236]^x[237]^x[238]^x[239]^x[240]^x[242]^x[243]^x[247]^x[251]^x[252]^x[253]^x[255]^x[257]^x[258]^x[259]^x[260]^x[262]^x[265]^x[271]^x[272]^x[273]^x[275]^x[276]^x[277]^x[278]^x[279]^x[280]^x[281]^x[282]^x[283]^x[285]^x[286]^x[287]^x[288]^x[290]^x[292]^x[293]^x[295]^x[298]^x[299]^u[63]^u[62]^u[61]^u[60]^u[59]^u[57]^u[56]^u[52]^u[48]^u[47]^u[46]^u[44]^u[42]^u[41]^u[40]^u[39]^u[37]^u[34]^u[28]^u[27]^u[26]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[14]^u[13]^u[12]^u[11]^u[9]^u[7]^u[6]^u[4]^u[1]^u[0];
	y[45] = x[236]^x[237]^x[240]^x[243]^x[244]^x[245]^x[248]^x[252]^x[253]^x[254]^x[255]^x[256]^x[258]^x[259]^x[261]^x[263]^x[264]^x[266]^x[269]^x[271]^x[272]^x[273]^x[274]^x[277]^x[278]^x[281]^x[282]^x[283]^x[284]^x[285]^x[286]^x[288]^x[291]^x[292]^x[295]^x[296]^x[298]^x[299]^u[63]^u[62]^u[59]^u[56]^u[55]^u[54]^u[51]^u[47]^u[46]^u[45]^u[44]^u[43]^u[41]^u[40]^u[38]^u[36]^u[35]^u[33]^u[30]^u[28]^u[27]^u[26]^u[25]^u[22]^u[21]^u[18]^u[17]^u[16]^u[15]^u[14]^u[13]^u[11]^u[8]^u[7]^u[4]^u[3]^u[1]^u[0];
	y[46] = x[236]^x[237]^x[239]^x[244]^x[246]^x[249]^x[253]^x[254]^x[256]^x[257]^x[259]^x[262]^x[265]^x[267]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[278]^x[280]^x[282]^x[283]^x[284]^x[286]^x[294]^x[295]^x[296]^x[297]^x[298]^x[299]^u[63]^u[62]^u[60]^u[55]^u[53]^u[50]^u[46]^u[45]^u[43]^u[42]^u[40]^u[37]^u[34]^u[32]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[21]^u[19]^u[17]^u[16]^u[15]^u[13]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[47] = x[236]^x[237]^x[239]^x[240]^x[241]^x[247]^x[250]^x[254]^x[257]^x[258]^x[263]^x[264]^x[266]^x[268]^x[269]^x[270]^x[272]^x[273]^x[274]^x[275]^x[277]^x[280]^x[281]^x[283]^x[284]^x[289]^x[292]^x[293]^x[294]^x[296]^x[297]^x[299]^u[63]^u[62]^u[60]^u[59]^u[58]^u[52]^u[49]^u[45]^u[42]^u[41]^u[36]^u[35]^u[33]^u[31]^u[30]^u[29]^u[27]^u[26]^u[25]^u[24]^u[22]^u[19]^u[18]^u[16]^u[15]^u[10]^u[7]^u[6]^u[5]^u[3]^u[2]^u[0];
	y[48] = x[236]^x[237]^x[239]^x[240]^x[242]^x[245]^x[248]^x[251]^x[258]^x[259]^x[260]^x[265]^x[267]^x[270]^x[273]^x[274]^x[275]^x[278]^x[279]^x[280]^x[281]^x[282]^x[284]^x[287]^x[289]^x[290]^x[292]^x[297]^u[63]^u[62]^u[60]^u[59]^u[57]^u[54]^u[51]^u[48]^u[41]^u[40]^u[39]^u[34]^u[32]^u[29]^u[26]^u[25]^u[24]^u[21]^u[20]^u[19]^u[18]^u[17]^u[15]^u[12]^u[10]^u[9]^u[7]^u[2];
	y[49] = x[237]^x[238]^x[240]^x[241]^x[243]^x[246]^x[249]^x[252]^x[259]^x[260]^x[261]^x[266]^x[268]^x[271]^x[274]^x[275]^x[276]^x[279]^x[280]^x[281]^x[282]^x[283]^x[285]^x[288]^x[290]^x[291]^x[293]^x[298]^u[62]^u[61]^u[59]^u[58]^u[56]^u[53]^u[50]^u[47]^u[40]^u[39]^u[38]^u[33]^u[31]^u[28]^u[25]^u[24]^u[23]^u[20]^u[19]^u[18]^u[17]^u[16]^u[14]^u[11]^u[9]^u[8]^u[6]^u[1];
	y[50] = x[236]^x[242]^x[244]^x[245]^x[247]^x[250]^x[253]^x[255]^x[261]^x[262]^x[264]^x[267]^x[271]^x[272]^x[275]^x[277]^x[279]^x[281]^x[282]^x[283]^x[284]^x[285]^x[286]^x[287]^x[291]^x[293]^x[295]^x[298]^x[299]^u[63]^u[57]^u[55]^u[54]^u[52]^u[49]^u[46]^u[44]^u[38]^u[37]^u[35]^u[32]^u[28]^u[27]^u[24]^u[22]^u[20]^u[18]^u[17]^u[16]^u[15]^u[14]^u[13]^u[12]^u[8]^u[6]^u[4]^u[1]^u[0];
	y[51] = x[236]^x[237]^x[238]^x[239]^x[241]^x[243]^x[246]^x[248]^x[251]^x[254]^x[255]^x[256]^x[260]^x[262]^x[263]^x[264]^x[265]^x[268]^x[269]^x[271]^x[272]^x[273]^x[278]^x[279]^x[282]^x[283]^x[284]^x[286]^x[288]^x[289]^x[293]^x[295]^x[296]^x[298]^x[299]^u[63]^u[62]^u[61]^u[60]^u[58]^u[56]^u[53]^u[51]^u[48]^u[45]^u[44]^u[43]^u[39]^u[37]^u[36]^u[35]^u[34]^u[31]^u[30]^u[28]^u[27]^u[26]^u[21]^u[20]^u[17]^u[16]^u[15]^u[13]^u[11]^u[10]^u[6]^u[4]^u[3]^u[1]^u[0];
	y[52] = x[236]^x[237]^x[240]^x[241]^x[242]^x[244]^x[245]^x[247]^x[249]^x[252]^x[256]^x[257]^x[260]^x[261]^x[263]^x[265]^x[266]^x[270]^x[271]^x[272]^x[273]^x[274]^x[276]^x[283]^x[284]^x[290]^x[292]^x[293]^x[295]^x[296]^x[297]^x[298]^x[299]^u[63]^u[62]^u[59]^u[58]^u[57]^u[55]^u[54]^u[52]^u[50]^u[47]^u[43]^u[42]^u[39]^u[38]^u[36]^u[34]^u[33]^u[29]^u[28]^u[27]^u[26]^u[25]^u[23]^u[16]^u[15]^u[9]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[53] = x[237]^x[238]^x[241]^x[242]^x[243]^x[245]^x[246]^x[248]^x[250]^x[253]^x[257]^x[258]^x[261]^x[262]^x[264]^x[266]^x[267]^x[271]^x[272]^x[273]^x[274]^x[275]^x[277]^x[284]^x[285]^x[291]^x[293]^x[294]^x[296]^x[297]^x[298]^x[299]^u[62]^u[61]^u[58]^u[57]^u[56]^u[54]^u[53]^u[51]^u[49]^u[46]^u[42]^u[41]^u[38]^u[37]^u[35]^u[33]^u[32]^u[28]^u[27]^u[26]^u[25]^u[24]^u[22]^u[15]^u[14]^u[8]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[54] = x[236]^x[241]^x[242]^x[243]^x[244]^x[245]^x[246]^x[247]^x[249]^x[251]^x[254]^x[255]^x[258]^x[259]^x[260]^x[262]^x[263]^x[264]^x[265]^x[267]^x[268]^x[269]^x[271]^x[272]^x[273]^x[274]^x[275]^x[278]^x[279]^x[280]^x[286]^x[287]^x[289]^x[293]^x[297]^x[299]^u[63]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[52]^u[50]^u[48]^u[45]^u[44]^u[41]^u[40]^u[39]^u[37]^u[36]^u[35]^u[34]^u[32]^u[31]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[21]^u[20]^u[19]^u[13]^u[12]^u[10]^u[6]^u[2]^u[0];
	y[55] = x[236]^x[237]^x[238]^x[239]^x[241]^x[242]^x[243]^x[244]^x[246]^x[247]^x[248]^x[250]^x[252]^x[256]^x[259]^x[261]^x[263]^x[265]^x[266]^x[268]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[281]^x[285]^x[288]^x[289]^x[290]^x[292]^x[293]^x[295]^u[63]^u[62]^u[61]^u[60]^u[58]^u[57]^u[56]^u[55]^u[53]^u[52]^u[51]^u[49]^u[47]^u[43]^u[40]^u[38]^u[36]^u[34]^u[33]^u[31]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[18]^u[14]^u[11]^u[10]^u[9]^u[7]^u[6]^u[4];
	y[56] = x[237]^x[238]^x[239]^x[240]^x[242]^x[243]^x[244]^x[245]^x[247]^x[248]^x[249]^x[251]^x[253]^x[257]^x[260]^x[262]^x[264]^x[266]^x[267]^x[269]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[282]^x[286]^x[289]^x[290]^x[291]^x[293]^x[294]^x[296]^u[62]^u[61]^u[60]^u[59]^u[57]^u[56]^u[55]^u[54]^u[52]^u[51]^u[50]^u[48]^u[46]^u[42]^u[39]^u[37]^u[35]^u[33]^u[32]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[17]^u[13]^u[10]^u[9]^u[8]^u[6]^u[5]^u[3];
	y[57] = x[236]^x[240]^x[243]^x[244]^x[246]^x[248]^x[249]^x[250]^x[252]^x[254]^x[255]^x[258]^x[260]^x[261]^x[263]^x[264]^x[265]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[277]^x[279]^x[280]^x[283]^x[285]^x[289]^x[290]^x[291]^x[293]^x[297]^x[298]^u[63]^u[59]^u[56]^u[55]^u[53]^u[51]^u[50]^u[49]^u[47]^u[45]^u[44]^u[41]^u[39]^u[38]^u[36]^u[35]^u[34]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[22]^u[20]^u[19]^u[16]^u[14]^u[10]^u[9]^u[8]^u[6]^u[2]^u[1];
	y[58] = x[237]^x[241]^x[244]^x[245]^x[247]^x[249]^x[250]^x[251]^x[253]^x[255]^x[256]^x[259]^x[261]^x[262]^x[264]^x[265]^x[266]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[278]^x[280]^x[281]^x[284]^x[286]^x[290]^x[291]^x[292]^x[294]^x[298]^x[299]^u[62]^u[58]^u[55]^u[54]^u[52]^u[50]^u[49]^u[48]^u[46]^u[44]^u[43]^u[40]^u[38]^u[37]^u[35]^u[34]^u[33]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[21]^u[19]^u[18]^u[15]^u[13]^u[9]^u[8]^u[7]^u[5]^u[1]^u[0];
	y[59] = x[238]^x[242]^x[245]^x[246]^x[248]^x[250]^x[251]^x[252]^x[254]^x[256]^x[257]^x[260]^x[262]^x[263]^x[265]^x[266]^x[267]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[277]^x[279]^x[281]^x[282]^x[285]^x[287]^x[291]^x[292]^x[293]^x[295]^x[299]^u[61]^u[57]^u[54]^u[53]^u[51]^u[49]^u[48]^u[47]^u[45]^u[43]^u[42]^u[39]^u[37]^u[36]^u[34]^u[33]^u[32]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[20]^u[18]^u[17]^u[14]^u[12]^u[8]^u[7]^u[6]^u[4]^u[0];
	y[60] = x[236]^x[238]^x[241]^x[243]^x[245]^x[246]^x[247]^x[249]^x[251]^x[252]^x[253]^x[257]^x[258]^x[260]^x[261]^x[263]^x[266]^x[267]^x[268]^x[269]^x[270]^x[272]^x[273]^x[274]^x[275]^x[277]^x[278]^x[279]^x[282]^x[283]^x[285]^x[286]^x[287]^x[288]^x[289]^x[295]^x[296]^x[298]^u[63]^u[61]^u[58]^u[56]^u[54]^u[53]^u[52]^u[50]^u[48]^u[47]^u[46]^u[42]^u[41]^u[39]^u[38]^u[36]^u[33]^u[32]^u[31]^u[30]^u[29]^u[27]^u[26]^u[25]^u[24]^u[22]^u[21]^u[20]^u[17]^u[16]^u[14]^u[13]^u[12]^u[11]^u[10]^u[4]^u[3]^u[1];
	y[61] = x[237]^x[239]^x[242]^x[244]^x[246]^x[247]^x[248]^x[250]^x[252]^x[253]^x[254]^x[258]^x[259]^x[261]^x[262]^x[264]^x[267]^x[268]^x[269]^x[270]^x[271]^x[273]^x[274]^x[275]^x[276]^x[278]^x[279]^x[280]^x[283]^x[284]^x[286]^x[287]^x[288]^x[289]^x[290]^x[296]^x[297]^x[299]^u[62]^u[60]^u[57]^u[55]^u[53]^u[52]^u[51]^u[49]^u[47]^u[46]^u[45]^u[41]^u[40]^u[38]^u[37]^u[35]^u[32]^u[31]^u[30]^u[29]^u[28]^u[26]^u[25]^u[24]^u[23]^u[21]^u[20]^u[19]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[9]^u[3]^u[2]^u[0];
	y[62] = x[236]^x[239]^x[240]^x[241]^x[243]^x[247]^x[248]^x[249]^x[251]^x[253]^x[254]^x[259]^x[262]^x[263]^x[264]^x[265]^x[268]^x[270]^x[272]^x[274]^x[275]^x[277]^x[281]^x[284]^x[288]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[297]^u[63]^u[60]^u[59]^u[58]^u[56]^u[52]^u[51]^u[50]^u[48]^u[46]^u[45]^u[40]^u[37]^u[36]^u[35]^u[34]^u[31]^u[29]^u[27]^u[25]^u[24]^u[22]^u[18]^u[15]^u[11]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[2];
	y[63] = x[236]^x[237]^x[238]^x[239]^x[240]^x[242]^x[244]^x[245]^x[248]^x[249]^x[250]^x[252]^x[254]^x[263]^x[265]^x[266]^x[273]^x[275]^x[278]^x[279]^x[280]^x[282]^x[287]^x[291]^x[296]^u[63]^u[62]^u[61]^u[60]^u[59]^u[57]^u[55]^u[54]^u[51]^u[50]^u[49]^u[47]^u[45]^u[36]^u[34]^u[33]^u[26]^u[24]^u[21]^u[20]^u[19]^u[17]^u[12]^u[8]^u[3];
	y[64] = x[0]^x[236]^x[237]^x[240]^x[243]^x[246]^x[249]^x[250]^x[251]^x[253]^x[260]^x[266]^x[267]^x[269]^x[271]^x[274]^x[281]^x[283]^x[285]^x[287]^x[288]^x[289]^x[293]^x[294]^x[295]^x[297]^x[298]^u[63]^u[62]^u[59]^u[56]^u[53]^u[50]^u[49]^u[48]^u[46]^u[39]^u[33]^u[32]^u[30]^u[28]^u[25]^u[18]^u[16]^u[14]^u[12]^u[11]^u[10]^u[6]^u[5]^u[4]^u[2]^u[1];
	y[65] = x[1]^x[236]^x[237]^x[239]^x[244]^x[245]^x[247]^x[250]^x[251]^x[252]^x[254]^x[255]^x[260]^x[261]^x[264]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[275]^x[276]^x[279]^x[280]^x[282]^x[284]^x[285]^x[286]^x[287]^x[288]^x[290]^x[292]^x[293]^x[296]^x[299]^u[63]^u[62]^u[60]^u[55]^u[54]^u[52]^u[49]^u[48]^u[47]^u[45]^u[44]^u[39]^u[38]^u[35]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[24]^u[23]^u[20]^u[19]^u[17]^u[15]^u[14]^u[13]^u[12]^u[11]^u[9]^u[7]^u[6]^u[3]^u[0];
	y[66] = x[2]^x[236]^x[237]^x[239]^x[240]^x[241]^x[246]^x[248]^x[251]^x[252]^x[253]^x[256]^x[260]^x[261]^x[262]^x[264]^x[265]^x[268]^x[270]^x[272]^x[273]^x[277]^x[279]^x[281]^x[283]^x[286]^x[288]^x[291]^x[292]^x[295]^x[297]^x[298]^u[63]^u[62]^u[60]^u[59]^u[58]^u[53]^u[51]^u[48]^u[47]^u[46]^u[43]^u[39]^u[38]^u[37]^u[35]^u[34]^u[31]^u[29]^u[27]^u[26]^u[22]^u[20]^u[18]^u[16]^u[13]^u[11]^u[8]^u[7]^u[4]^u[2]^u[1];
	y[67] = x[3]^x[236]^x[237]^x[239]^x[240]^x[242]^x[245]^x[247]^x[249]^x[252]^x[253]^x[254]^x[255]^x[257]^x[260]^x[261]^x[262]^x[263]^x[264]^x[265]^x[266]^x[273]^x[274]^x[276]^x[278]^x[279]^x[282]^x[284]^x[285]^x[294]^x[295]^x[296]^x[299]^u[63]^u[62]^u[60]^u[59]^u[57]^u[54]^u[52]^u[50]^u[47]^u[46]^u[45]^u[44]^u[42]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[26]^u[25]^u[23]^u[21]^u[20]^u[17]^u[15]^u[14]^u[5]^u[4]^u[3]^u[0];
	y[68] = x[4]^x[236]^x[237]^x[239]^x[240]^x[243]^x[245]^x[246]^x[248]^x[250]^x[253]^x[254]^x[256]^x[258]^x[260]^x[261]^x[262]^x[263]^x[265]^x[266]^x[267]^x[269]^x[271]^x[274]^x[275]^x[276]^x[277]^x[283]^x[286]^x[287]^x[289]^x[292]^x[293]^x[294]^x[296]^x[297]^x[298]^u[63]^u[62]^u[60]^u[59]^u[56]^u[54]^u[53]^u[51]^u[49]^u[46]^u[45]^u[43]^u[41]^u[39]^u[38]^u[37]^u[36]^u[34]^u[33]^u[32]^u[30]^u[28]^u[25]^u[24]^u[23]^u[22]^u[16]^u[13]^u[12]^u[10]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[69] = x[5]^x[237]^x[238]^x[240]^x[241]^x[244]^x[246]^x[247]^x[249]^x[251]^x[254]^x[255]^x[257]^x[259]^x[261]^x[262]^x[263]^x[264]^x[266]^x[267]^x[268]^x[270]^x[272]^x[275]^x[276]^x[277]^x[278]^x[284]^x[287]^x[288]^x[290]^x[293]^x[294]^x[295]^x[297]^x[298]^x[299]^u[62]^u[61]^u[59]^u[58]^u[55]^u[53]^u[52]^u[50]^u[48]^u[45]^u[44]^u[42]^u[40]^u[38]^u[37]^u[36]^u[35]^u[33]^u[32]^u[31]^u[29]^u[27]^u[24]^u[23]^u[22]^u[21]^u[15]^u[12]^u[11]^u[9]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[70] = x[6]^x[238]^x[239]^x[241]^x[242]^x[245]^x[247]^x[248]^x[250]^x[252]^x[255]^x[256]^x[258]^x[260]^x[262]^x[263]^x[264]^x[265]^x[267]^x[268]^x[269]^x[271]^x[273]^x[276]^x[277]^x[278]^x[279]^x[285]^x[288]^x[289]^x[291]^x[294]^x[295]^x[296]^x[298]^x[299]^u[61]^u[60]^u[58]^u[57]^u[54]^u[52]^u[51]^u[49]^u[47]^u[44]^u[43]^u[41]^u[39]^u[37]^u[36]^u[35]^u[34]^u[32]^u[31]^u[30]^u[28]^u[26]^u[23]^u[22]^u[21]^u[20]^u[14]^u[11]^u[10]^u[8]^u[5]^u[4]^u[3]^u[1]^u[0];
	y[71] = x[7]^x[239]^x[240]^x[242]^x[243]^x[246]^x[248]^x[249]^x[251]^x[253]^x[256]^x[257]^x[259]^x[261]^x[263]^x[264]^x[265]^x[266]^x[268]^x[269]^x[270]^x[272]^x[274]^x[277]^x[278]^x[279]^x[280]^x[286]^x[289]^x[290]^x[292]^x[295]^x[296]^x[297]^x[299]^u[60]^u[59]^u[57]^u[56]^u[53]^u[51]^u[50]^u[48]^u[46]^u[43]^u[42]^u[40]^u[38]^u[36]^u[35]^u[34]^u[33]^u[31]^u[30]^u[29]^u[27]^u[25]^u[22]^u[21]^u[20]^u[19]^u[13]^u[10]^u[9]^u[7]^u[4]^u[3]^u[2]^u[0];
	y[72] = x[8]^x[240]^x[241]^x[243]^x[244]^x[247]^x[249]^x[250]^x[252]^x[254]^x[257]^x[258]^x[260]^x[262]^x[264]^x[265]^x[266]^x[267]^x[269]^x[270]^x[271]^x[273]^x[275]^x[278]^x[279]^x[280]^x[281]^x[287]^x[290]^x[291]^x[293]^x[296]^x[297]^x[298]^u[59]^u[58]^u[56]^u[55]^u[52]^u[50]^u[49]^u[47]^u[45]^u[42]^u[41]^u[39]^u[37]^u[35]^u[34]^u[33]^u[32]^u[30]^u[29]^u[28]^u[26]^u[24]^u[21]^u[20]^u[19]^u[18]^u[12]^u[9]^u[8]^u[6]^u[3]^u[2]^u[1];
	y[73] = x[9]^x[236]^x[238]^x[239]^x[242]^x[244]^x[248]^x[250]^x[251]^x[253]^x[258]^x[259]^x[260]^x[261]^x[263]^x[264]^x[265]^x[266]^x[267]^x[268]^x[269]^x[270]^x[272]^x[274]^x[281]^x[282]^x[285]^x[287]^x[288]^x[289]^x[291]^x[293]^x[295]^x[297]^x[299]^u[63]^u[61]^u[60]^u[57]^u[55]^u[51]^u[49]^u[48]^u[46]^u[41]^u[40]^u[39]^u[38]^u[36]^u[35]^u[34]^u[33]^u[32]^u[31]^u[30]^u[29]^u[27]^u[25]^u[18]^u[17]^u[14]^u[12]^u[11]^u[10]^u[8]^u[6]^u[4]^u[2]^u[0];
	y[74] = x[10]^x[236]^x[237]^x[238]^x[240]^x[241]^x[243]^x[249]^x[251]^x[252]^x[254]^x[255]^x[259]^x[261]^x[262]^x[265]^x[266]^x[267]^x[268]^x[270]^x[273]^x[275]^x[276]^x[279]^x[280]^x[282]^x[283]^x[285]^x[286]^x[287]^x[288]^x[290]^x[293]^x[295]^x[296]^u[63]^u[62]^u[61]^u[59]^u[58]^u[56]^u[50]^u[48]^u[47]^u[45]^u[44]^u[40]^u[38]^u[37]^u[34]^u[33]^u[32]^u[31]^u[29]^u[26]^u[24]^u[23]^u[20]^u[19]^u[17]^u[16]^u[14]^u[13]^u[12]^u[11]^u[9]^u[6]^u[4]^u[3];
	y[75] = x[11]^x[236]^x[237]^x[242]^x[244]^x[245]^x[250]^x[252]^x[253]^x[256]^x[262]^x[263]^x[264]^x[266]^x[267]^x[268]^x[274]^x[277]^x[279]^x[281]^x[283]^x[284]^x[285]^x[286]^x[288]^x[291]^x[292]^x[293]^x[295]^x[296]^x[297]^x[298]^u[63]^u[62]^u[57]^u[55]^u[54]^u[49]^u[47]^u[46]^u[43]^u[37]^u[36]^u[35]^u[33]^u[32]^u[31]^u[25]^u[22]^u[20]^u[18]^u[16]^u[15]^u[14]^u[13]^u[11]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1];
	y[76] = x[12]^x[237]^x[238]^x[243]^x[245]^x[246]^x[251]^x[253]^x[254]^x[257]^x[263]^x[264]^x[265]^x[267]^x[268]^x[269]^x[275]^x[278]^x[280]^x[282]^x[284]^x[285]^x[286]^x[287]^x[289]^x[292]^x[293]^x[294]^x[296]^x[297]^x[298]^x[299]^u[62]^u[61]^u[56]^u[54]^u[53]^u[48]^u[46]^u[45]^u[42]^u[36]^u[35]^u[34]^u[32]^u[31]^u[30]^u[24]^u[21]^u[19]^u[17]^u[15]^u[14]^u[13]^u[12]^u[10]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[77] = x[13]^x[238]^x[239]^x[244]^x[246]^x[247]^x[252]^x[254]^x[255]^x[258]^x[264]^x[265]^x[266]^x[268]^x[269]^x[270]^x[276]^x[279]^x[281]^x[283]^x[285]^x[286]^x[287]^x[288]^x[290]^x[293]^x[294]^x[295]^x[297]^x[298]^x[299]^u[61]^u[60]^u[55]^u[53]^u[52]^u[47]^u[45]^u[44]^u[41]^u[35]^u[34]^u[33]^u[31]^u[30]^u[29]^u[23]^u[20]^u[18]^u[16]^u[14]^u[13]^u[12]^u[11]^u[9]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[78] = x[14]^x[236]^x[238]^x[240]^x[241]^x[247]^x[248]^x[253]^x[256]^x[259]^x[260]^x[264]^x[265]^x[266]^x[267]^x[270]^x[276]^x[277]^x[279]^x[282]^x[284]^x[285]^x[286]^x[288]^x[291]^x[292]^x[293]^x[296]^x[299]^u[63]^u[61]^u[59]^u[58]^u[52]^u[51]^u[46]^u[43]^u[40]^u[39]^u[35]^u[34]^u[33]^u[32]^u[29]^u[23]^u[22]^u[20]^u[17]^u[15]^u[14]^u[13]^u[11]^u[8]^u[7]^u[6]^u[3]^u[0];
	y[79] = x[15]^x[237]^x[239]^x[241]^x[242]^x[248]^x[249]^x[254]^x[257]^x[260]^x[261]^x[265]^x[266]^x[267]^x[268]^x[271]^x[277]^x[278]^x[280]^x[283]^x[285]^x[286]^x[287]^x[289]^x[292]^x[293]^x[294]^x[297]^u[62]^u[60]^u[58]^u[57]^u[51]^u[50]^u[45]^u[42]^u[39]^u[38]^u[34]^u[33]^u[32]^u[31]^u[28]^u[22]^u[21]^u[19]^u[16]^u[14]^u[13]^u[12]^u[10]^u[7]^u[6]^u[5]^u[2];
	y[80] = x[16]^x[238]^x[240]^x[242]^x[243]^x[249]^x[250]^x[255]^x[258]^x[261]^x[262]^x[266]^x[267]^x[268]^x[269]^x[272]^x[278]^x[279]^x[281]^x[284]^x[286]^x[287]^x[288]^x[290]^x[293]^x[294]^x[295]^x[298]^u[61]^u[59]^u[57]^u[56]^u[50]^u[49]^u[44]^u[41]^u[38]^u[37]^u[33]^u[32]^u[31]^u[30]^u[27]^u[21]^u[20]^u[18]^u[15]^u[13]^u[12]^u[11]^u[9]^u[6]^u[5]^u[4]^u[1];
	y[81] = x[17]^x[236]^x[238]^x[243]^x[244]^x[245]^x[250]^x[251]^x[255]^x[256]^x[259]^x[260]^x[262]^x[263]^x[264]^x[267]^x[268]^x[270]^x[271]^x[273]^x[276]^x[282]^x[288]^x[291]^x[292]^x[293]^x[296]^x[298]^x[299]^u[63]^u[61]^u[56]^u[55]^u[54]^u[49]^u[48]^u[44]^u[43]^u[40]^u[39]^u[37]^u[36]^u[35]^u[32]^u[31]^u[29]^u[28]^u[26]^u[23]^u[17]^u[11]^u[8]^u[7]^u[6]^u[3]^u[1]^u[0];
	y[82] = x[18]^x[237]^x[239]^x[244]^x[245]^x[246]^x[251]^x[252]^x[256]^x[257]^x[260]^x[261]^x[263]^x[264]^x[265]^x[268]^x[269]^x[271]^x[272]^x[274]^x[277]^x[283]^x[289]^x[292]^x[293]^x[294]^x[297]^x[299]^u[62]^u[60]^u[55]^u[54]^u[53]^u[48]^u[47]^u[43]^u[42]^u[39]^u[38]^u[36]^u[35]^u[34]^u[31]^u[30]^u[28]^u[27]^u[25]^u[22]^u[16]^u[10]^u[7]^u[6]^u[5]^u[2]^u[0];
	y[83] = x[19]^x[238]^x[240]^x[245]^x[246]^x[247]^x[252]^x[253]^x[257]^x[258]^x[261]^x[262]^x[264]^x[265]^x[266]^x[269]^x[270]^x[272]^x[273]^x[275]^x[278]^x[284]^x[290]^x[293]^x[294]^x[295]^x[298]^u[61]^u[59]^u[54]^u[53]^u[52]^u[47]^u[46]^u[42]^u[41]^u[38]^u[37]^u[35]^u[34]^u[33]^u[30]^u[29]^u[27]^u[26]^u[24]^u[21]^u[15]^u[9]^u[6]^u[5]^u[4]^u[1];
	y[84] = x[20]^x[239]^x[241]^x[246]^x[247]^x[248]^x[253]^x[254]^x[258]^x[259]^x[262]^x[263]^x[265]^x[266]^x[267]^x[270]^x[271]^x[273]^x[274]^x[276]^x[279]^x[285]^x[291]^x[294]^x[295]^x[296]^x[299]^u[60]^u[58]^u[53]^u[52]^u[51]^u[46]^u[45]^u[41]^u[40]^u[37]^u[36]^u[34]^u[33]^u[32]^u[29]^u[28]^u[26]^u[25]^u[23]^u[20]^u[14]^u[8]^u[5]^u[4]^u[3]^u[0];
	y[85] = x[21]^x[240]^x[242]^x[247]^x[248]^x[249]^x[254]^x[255]^x[259]^x[260]^x[263]^x[264]^x[266]^x[267]^x[268]^x[271]^x[272]^x[274]^x[275]^x[277]^x[280]^x[286]^x[292]^x[295]^x[296]^x[297]^u[59]^u[57]^u[52]^u[51]^u[50]^u[45]^u[44]^u[40]^u[39]^u[36]^u[35]^u[33]^u[32]^u[31]^u[28]^u[27]^u[25]^u[24]^u[22]^u[19]^u[13]^u[7]^u[4]^u[3]^u[2];
	y[86] = x[22]^x[236]^x[238]^x[239]^x[243]^x[245]^x[248]^x[249]^x[250]^x[256]^x[261]^x[265]^x[267]^x[268]^x[271]^x[272]^x[273]^x[275]^x[278]^x[279]^x[280]^x[281]^x[285]^x[289]^x[292]^x[294]^x[295]^x[296]^x[297]^u[63]^u[61]^u[60]^u[56]^u[54]^u[51]^u[50]^u[49]^u[43]^u[38]^u[34]^u[32]^u[31]^u[28]^u[27]^u[26]^u[24]^u[21]^u[20]^u[19]^u[18]^u[14]^u[10]^u[7]^u[5]^u[4]^u[3]^u[2];
	y[87] = x[23]^x[237]^x[239]^x[240]^x[244]^x[246]^x[249]^x[250]^x[251]^x[257]^x[262]^x[266]^x[268]^x[269]^x[272]^x[273]^x[274]^x[276]^x[279]^x[280]^x[281]^x[282]^x[286]^x[290]^x[293]^x[295]^x[296]^x[297]^x[298]^u[62]^u[60]^u[59]^u[55]^u[53]^u[50]^u[49]^u[48]^u[42]^u[37]^u[33]^u[31]^u[30]^u[27]^u[26]^u[25]^u[23]^u[20]^u[19]^u[18]^u[17]^u[13]^u[9]^u[6]^u[4]^u[3]^u[2]^u[1];
	y[88] = x[24]^x[236]^x[239]^x[240]^x[247]^x[250]^x[251]^x[252]^x[255]^x[258]^x[260]^x[263]^x[264]^x[267]^x[270]^x[271]^x[273]^x[274]^x[275]^x[276]^x[277]^x[279]^x[281]^x[282]^x[283]^x[285]^x[289]^x[291]^x[292]^x[293]^x[295]^x[296]^x[297]^x[299]^u[63]^u[60]^u[59]^u[52]^u[49]^u[48]^u[47]^u[44]^u[41]^u[39]^u[36]^u[35]^u[32]^u[29]^u[28]^u[26]^u[25]^u[24]^u[23]^u[22]^u[20]^u[18]^u[17]^u[16]^u[14]^u[10]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[0];
	y[89] = x[25]^x[237]^x[240]^x[241]^x[248]^x[251]^x[252]^x[253]^x[256]^x[259]^x[261]^x[264]^x[265]^x[268]^x[271]^x[272]^x[274]^x[275]^x[276]^x[277]^x[278]^x[280]^x[282]^x[283]^x[284]^x[286]^x[290]^x[292]^x[293]^x[294]^x[296]^x[297]^x[298]^u[62]^u[59]^u[58]^u[51]^u[48]^u[47]^u[46]^u[43]^u[40]^u[38]^u[35]^u[34]^u[31]^u[28]^u[27]^u[25]^u[24]^u[23]^u[22]^u[21]^u[19]^u[17]^u[16]^u[15]^u[13]^u[9]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[90] = x[26]^x[236]^x[239]^x[242]^x[245]^x[249]^x[252]^x[253]^x[254]^x[255]^x[257]^x[262]^x[264]^x[265]^x[266]^x[271]^x[272]^x[273]^x[275]^x[277]^x[278]^x[280]^x[281]^x[283]^x[284]^x[289]^x[291]^x[292]^x[297]^x[299]^u[63]^u[60]^u[57]^u[54]^u[50]^u[47]^u[46]^u[45]^u[44]^u[42]^u[37]^u[35]^u[34]^u[33]^u[28]^u[27]^u[26]^u[24]^u[22]^u[21]^u[19]^u[18]^u[16]^u[15]^u[10]^u[8]^u[7]^u[2]^u[0];
	y[91] = x[27]^x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[243]^x[245]^x[246]^x[250]^x[253]^x[254]^x[256]^x[258]^x[260]^x[263]^x[264]^x[265]^x[266]^x[267]^x[269]^x[271]^x[272]^x[273]^x[274]^x[278]^x[280]^x[281]^x[282]^x[284]^x[287]^x[289]^x[290]^x[294]^x[295]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[56]^u[54]^u[53]^u[49]^u[46]^u[45]^u[43]^u[41]^u[39]^u[36]^u[35]^u[34]^u[33]^u[32]^u[30]^u[28]^u[27]^u[26]^u[25]^u[21]^u[19]^u[18]^u[17]^u[15]^u[12]^u[10]^u[9]^u[5]^u[4];
	y[92] = x[28]^x[236]^x[237]^x[240]^x[242]^x[244]^x[245]^x[246]^x[247]^x[251]^x[254]^x[257]^x[259]^x[260]^x[261]^x[265]^x[266]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[280]^x[281]^x[282]^x[283]^x[287]^x[288]^x[289]^x[290]^x[291]^x[292]^x[293]^x[294]^x[296]^x[298]^u[63]^u[62]^u[59]^u[57]^u[55]^u[54]^u[53]^u[52]^u[48]^u[45]^u[42]^u[40]^u[39]^u[38]^u[34]^u[33]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[19]^u[18]^u[17]^u[16]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[3]^u[1];
	y[93] = x[29]^x[237]^x[238]^x[241]^x[243]^x[245]^x[246]^x[247]^x[248]^x[252]^x[255]^x[258]^x[260]^x[261]^x[262]^x[266]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[277]^x[281]^x[282]^x[283]^x[284]^x[288]^x[289]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[297]^x[299]^u[62]^u[61]^u[58]^u[56]^u[54]^u[53]^u[52]^u[51]^u[47]^u[44]^u[41]^u[39]^u[38]^u[37]^u[33]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[18]^u[17]^u[16]^u[15]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[2]^u[0];
	y[94] = x[30]^x[238]^x[239]^x[242]^x[244]^x[246]^x[247]^x[248]^x[249]^x[253]^x[256]^x[259]^x[261]^x[262]^x[263]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[277]^x[278]^x[282]^x[283]^x[284]^x[285]^x[289]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[296]^x[298]^u[61]^u[60]^u[57]^u[55]^u[53]^u[52]^u[51]^u[50]^u[46]^u[43]^u[40]^u[38]^u[37]^u[36]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[17]^u[16]^u[15]^u[14]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3]^u[1];
	y[95] = x[31]^x[239]^x[240]^x[243]^x[245]^x[247]^x[248]^x[249]^x[250]^x[254]^x[257]^x[260]^x[262]^x[263]^x[264]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[277]^x[278]^x[279]^x[283]^x[284]^x[285]^x[286]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[296]^x[297]^x[299]^u[60]^u[59]^u[56]^u[54]^u[52]^u[51]^u[50]^u[49]^u[45]^u[42]^u[39]^u[37]^u[36]^u[35]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[16]^u[15]^u[14]^u[13]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2]^u[0];
	y[96] = x[32]^x[240]^x[241]^x[244]^x[246]^x[248]^x[249]^x[250]^x[251]^x[255]^x[258]^x[261]^x[263]^x[264]^x[265]^x[269]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[277]^x[278]^x[279]^x[280]^x[284]^x[285]^x[286]^x[287]^x[291]^x[292]^x[293]^x[294]^x[295]^x[296]^x[297]^x[298]^u[59]^u[58]^u[55]^u[53]^u[51]^u[50]^u[49]^u[48]^u[44]^u[41]^u[38]^u[36]^u[35]^u[34]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[15]^u[14]^u[13]^u[12]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[97] = x[33]^x[236]^x[238]^x[239]^x[242]^x[247]^x[249]^x[250]^x[251]^x[252]^x[255]^x[256]^x[259]^x[260]^x[262]^x[265]^x[266]^x[269]^x[270]^x[272]^x[273]^x[274]^x[275]^x[277]^x[278]^x[281]^x[286]^x[288]^x[289]^x[296]^x[297]^x[299]^u[63]^u[61]^u[60]^u[57]^u[52]^u[50]^u[49]^u[48]^u[47]^u[44]^u[43]^u[40]^u[39]^u[37]^u[34]^u[33]^u[30]^u[29]^u[27]^u[26]^u[25]^u[24]^u[22]^u[21]^u[18]^u[13]^u[11]^u[10]^u[3]^u[2]^u[0];
	y[98] = x[34]^x[237]^x[239]^x[240]^x[243]^x[248]^x[250]^x[251]^x[252]^x[253]^x[256]^x[257]^x[260]^x[261]^x[263]^x[266]^x[267]^x[270]^x[271]^x[273]^x[274]^x[275]^x[276]^x[278]^x[279]^x[282]^x[287]^x[289]^x[290]^x[297]^x[298]^u[62]^u[60]^u[59]^u[56]^u[51]^u[49]^u[48]^u[47]^u[46]^u[43]^u[42]^u[39]^u[38]^u[36]^u[33]^u[32]^u[29]^u[28]^u[26]^u[25]^u[24]^u[23]^u[21]^u[20]^u[17]^u[12]^u[10]^u[9]^u[2]^u[1];
	y[99] = x[35]^x[236]^x[239]^x[240]^x[244]^x[245]^x[249]^x[251]^x[252]^x[253]^x[254]^x[255]^x[257]^x[258]^x[260]^x[261]^x[262]^x[267]^x[268]^x[269]^x[272]^x[274]^x[275]^x[277]^x[283]^x[285]^x[287]^x[288]^x[289]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[299]^u[63]^u[60]^u[59]^u[55]^u[54]^u[50]^u[48]^u[47]^u[46]^u[45]^u[44]^u[42]^u[41]^u[39]^u[38]^u[37]^u[32]^u[31]^u[30]^u[27]^u[25]^u[24]^u[22]^u[16]^u[14]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[0];
	y[100] = x[36]^x[237]^x[240]^x[241]^x[245]^x[246]^x[250]^x[252]^x[253]^x[254]^x[255]^x[256]^x[258]^x[259]^x[261]^x[262]^x[263]^x[268]^x[269]^x[270]^x[273]^x[275]^x[276]^x[278]^x[284]^x[286]^x[288]^x[289]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[296]^u[62]^u[59]^u[58]^u[54]^u[53]^u[49]^u[47]^u[46]^u[45]^u[44]^u[43]^u[41]^u[40]^u[38]^u[37]^u[36]^u[31]^u[30]^u[29]^u[26]^u[24]^u[23]^u[21]^u[15]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3];
	y[101] = x[37]^x[238]^x[241]^x[242]^x[246]^x[247]^x[251]^x[253]^x[254]^x[255]^x[256]^x[257]^x[259]^x[260]^x[262]^x[263]^x[264]^x[269]^x[270]^x[271]^x[274]^x[276]^x[277]^x[279]^x[285]^x[287]^x[289]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[296]^x[297]^u[61]^u[58]^u[57]^u[53]^u[52]^u[48]^u[46]^u[45]^u[44]^u[43]^u[42]^u[40]^u[39]^u[37]^u[36]^u[35]^u[30]^u[29]^u[28]^u[25]^u[23]^u[22]^u[20]^u[14]^u[12]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2];
	y[102] = x[38]^x[236]^x[238]^x[241]^x[242]^x[243]^x[245]^x[247]^x[248]^x[252]^x[254]^x[256]^x[257]^x[258]^x[261]^x[263]^x[265]^x[269]^x[270]^x[272]^x[275]^x[276]^x[277]^x[278]^x[279]^x[285]^x[286]^x[287]^x[288]^x[289]^x[290]^x[291]^x[296]^x[297]^u[63]^u[61]^u[58]^u[57]^u[56]^u[54]^u[52]^u[51]^u[47]^u[45]^u[43]^u[42]^u[41]^u[38]^u[36]^u[34]^u[30]^u[29]^u[27]^u[24]^u[23]^u[22]^u[21]^u[20]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[3]^u[2];
	y[103] = x[39]^x[236]^x[237]^x[238]^x[241]^x[242]^x[243]^x[244]^x[245]^x[246]^x[248]^x[249]^x[253]^x[257]^x[258]^x[259]^x[260]^x[262]^x[266]^x[269]^x[270]^x[273]^x[277]^x[278]^x[285]^x[286]^x[288]^x[290]^x[291]^x[293]^x[294]^x[295]^x[297]^u[63]^u[62]^u[61]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[51]^u[50]^u[46]^u[42]^u[41]^u[40]^u[39]^u[37]^u[33]^u[30]^u[29]^u[26]^u[22]^u[21]^u[14]^u[13]^u[11]^u[9]^u[8]^u[6]^u[5]^u[4]^u[2];
	y[104] = x[40]^x[236]^x[237]^x[241]^x[242]^x[243]^x[244]^x[246]^x[247]^x[249]^x[250]^x[254]^x[255]^x[258]^x[259]^x[261]^x[263]^x[264]^x[267]^x[269]^x[270]^x[274]^x[276]^x[278]^x[280]^x[285]^x[286]^x[291]^x[293]^x[296]^u[63]^u[62]^u[58]^u[57]^u[56]^u[55]^u[53]^u[52]^u[50]^u[49]^u[45]^u[44]^u[41]^u[40]^u[38]^u[36]^u[35]^u[32]^u[30]^u[29]^u[25]^u[23]^u[21]^u[19]^u[14]^u[13]^u[8]^u[6]^u[3];
	y[105] = x[41]^x[236]^x[237]^x[239]^x[241]^x[242]^x[243]^x[244]^x[247]^x[248]^x[250]^x[251]^x[256]^x[259]^x[262]^x[265]^x[268]^x[269]^x[270]^x[275]^x[276]^x[277]^x[280]^x[281]^x[285]^x[286]^x[289]^x[293]^x[295]^x[297]^x[298]^u[63]^u[62]^u[60]^u[58]^u[57]^u[56]^u[55]^u[52]^u[51]^u[49]^u[48]^u[43]^u[40]^u[37]^u[34]^u[31]^u[30]^u[29]^u[24]^u[23]^u[22]^u[19]^u[18]^u[14]^u[13]^u[10]^u[6]^u[4]^u[2]^u[1];
	y[106] = x[42]^x[236]^x[237]^x[239]^x[240]^x[241]^x[242]^x[243]^x[244]^x[248]^x[249]^x[251]^x[252]^x[255]^x[257]^x[263]^x[264]^x[266]^x[270]^x[277]^x[278]^x[279]^x[280]^x[281]^x[282]^x[285]^x[286]^x[289]^x[290]^x[292]^x[293]^x[295]^x[296]^x[299]^u[63]^u[62]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[51]^u[50]^u[48]^u[47]^u[44]^u[42]^u[36]^u[35]^u[33]^u[29]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[14]^u[13]^u[10]^u[9]^u[7]^u[6]^u[4]^u[3]^u[0];
	y[107] = x[43]^x[237]^x[238]^x[240]^x[241]^x[242]^x[243]^x[244]^x[245]^x[249]^x[250]^x[252]^x[253]^x[256]^x[258]^x[264]^x[265]^x[267]^x[271]^x[278]^x[279]^x[280]^x[281]^x[282]^x[283]^x[286]^x[287]^x[290]^x[291]^x[293]^x[294]^x[296]^x[297]^u[62]^u[61]^u[59]^u[58]^u[57]^u[56]^u[55]^u[54]^u[50]^u[49]^u[47]^u[46]^u[43]^u[41]^u[35]^u[34]^u[32]^u[28]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[13]^u[12]^u[9]^u[8]^u[6]^u[5]^u[3]^u[2];
	y[108] = x[44]^x[238]^x[239]^x[241]^x[242]^x[243]^x[244]^x[245]^x[246]^x[250]^x[251]^x[253]^x[254]^x[257]^x[259]^x[265]^x[266]^x[268]^x[272]^x[279]^x[280]^x[281]^x[282]^x[283]^x[284]^x[287]^x[288]^x[291]^x[292]^x[294]^x[295]^x[297]^x[298]^u[61]^u[60]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[49]^u[48]^u[46]^u[45]^u[42]^u[40]^u[34]^u[33]^u[31]^u[27]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[12]^u[11]^u[8]^u[7]^u[5]^u[4]^u[2]^u[1];
	y[109] = x[45]^x[236]^x[238]^x[240]^x[241]^x[242]^x[243]^x[244]^x[246]^x[247]^x[251]^x[252]^x[254]^x[258]^x[264]^x[266]^x[267]^x[271]^x[273]^x[276]^x[279]^x[281]^x[282]^x[283]^x[284]^x[287]^x[288]^x[294]^x[296]^x[299]^u[63]^u[61]^u[59]^u[58]^u[57]^u[56]^u[55]^u[53]^u[52]^u[48]^u[47]^u[45]^u[41]^u[35]^u[33]^u[32]^u[28]^u[26]^u[23]^u[20]^u[18]^u[17]^u[16]^u[15]^u[12]^u[11]^u[5]^u[3]^u[0];
	y[110] = x[46]^x[237]^x[239]^x[241]^x[242]^x[243]^x[244]^x[245]^x[247]^x[248]^x[252]^x[253]^x[255]^x[259]^x[265]^x[267]^x[268]^x[272]^x[274]^x[277]^x[280]^x[282]^x[283]^x[284]^x[285]^x[288]^x[289]^x[295]^x[297]^u[62]^u[60]^u[58]^u[57]^u[56]^u[55]^u[54]^u[52]^u[51]^u[47]^u[46]^u[44]^u[40]^u[34]^u[32]^u[31]^u[27]^u[25]^u[22]^u[19]^u[17]^u[16]^u[15]^u[14]^u[11]^u[10]^u[4]^u[2];
	y[111] = x[47]^x[236]^x[239]^x[240]^x[241]^x[242]^x[243]^x[244]^x[246]^x[248]^x[249]^x[253]^x[254]^x[255]^x[256]^x[264]^x[266]^x[268]^x[271]^x[273]^x[275]^x[276]^x[278]^x[279]^x[280]^x[281]^x[283]^x[284]^x[286]^x[287]^x[290]^x[292]^x[293]^x[294]^x[295]^x[296]^u[63]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[53]^u[51]^u[50]^u[46]^u[45]^u[44]^u[43]^u[35]^u[33]^u[31]^u[28]^u[26]^u[24]^u[23]^u[21]^u[20]^u[19]^u[18]^u[16]^u[15]^u[13]^u[12]^u[9]^u[7]^u[6]^u[5]^u[4]^u[3];
	y[112] = x[48]^x[236]^x[237]^x[238]^x[239]^x[240]^x[242]^x[243]^x[244]^x[247]^x[249]^x[250]^x[254]^x[256]^x[257]^x[260]^x[264]^x[265]^x[267]^x[271]^x[272]^x[274]^x[277]^x[281]^x[282]^x[284]^x[288]^x[289]^x[291]^x[292]^x[296]^x[297]^x[298]^u[63]^u[62]^u[61]^u[60]^u[59]^u[57]^u[56]^u[55]^u[52]^u[50]^u[49]^u[45]^u[43]^u[42]^u[39]^u[35]^u[34]^u[32]^u[28]^u[27]^u[25]^u[22]^u[18]^u[17]^u[15]^u[11]^u[10]^u[8]^u[7]^u[3]^u[2]^u[1];
	y[113] = x[49]^x[237]^x[238]^x[239]^x[240]^x[241]^x[243]^x[244]^x[245]^x[248]^x[250]^x[251]^x[255]^x[257]^x[258]^x[261]^x[265]^x[266]^x[268]^x[272]^x[273]^x[275]^x[278]^x[282]^x[283]^x[285]^x[289]^x[290]^x[292]^x[293]^x[297]^x[298]^x[299]^u[62]^u[61]^u[60]^u[59]^u[58]^u[56]^u[55]^u[54]^u[51]^u[49]^u[48]^u[44]^u[42]^u[41]^u[38]^u[34]^u[33]^u[31]^u[27]^u[26]^u[24]^u[21]^u[17]^u[16]^u[14]^u[10]^u[9]^u[7]^u[6]^u[2]^u[1]^u[0];
	y[114] = x[50]^x[236]^x[240]^x[242]^x[244]^x[246]^x[249]^x[251]^x[252]^x[255]^x[256]^x[258]^x[259]^x[260]^x[262]^x[264]^x[266]^x[267]^x[271]^x[273]^x[274]^x[280]^x[283]^x[284]^x[285]^x[286]^x[287]^x[289]^x[290]^x[291]^x[292]^x[295]^x[299]^u[63]^u[59]^u[57]^u[55]^u[53]^u[50]^u[48]^u[47]^u[44]^u[43]^u[41]^u[40]^u[39]^u[37]^u[35]^u[33]^u[32]^u[28]^u[26]^u[25]^u[19]^u[16]^u[15]^u[14]^u[13]^u[12]^u[10]^u[9]^u[8]^u[7]^u[4]^u[0];
	y[115] = x[51]^x[237]^x[241]^x[243]^x[245]^x[247]^x[250]^x[252]^x[253]^x[256]^x[257]^x[259]^x[260]^x[261]^x[263]^x[265]^x[267]^x[268]^x[272]^x[274]^x[275]^x[281]^x[284]^x[285]^x[286]^x[287]^x[288]^x[290]^x[291]^x[292]^x[293]^x[296]^u[62]^u[58]^u[56]^u[54]^u[52]^u[49]^u[47]^u[46]^u[43]^u[42]^u[40]^u[39]^u[38]^u[36]^u[34]^u[32]^u[31]^u[27]^u[25]^u[24]^u[18]^u[15]^u[14]^u[13]^u[12]^u[11]^u[9]^u[8]^u[7]^u[6]^u[3];
	y[116] = x[52]^x[238]^x[242]^x[244]^x[246]^x[248]^x[251]^x[253]^x[254]^x[257]^x[258]^x[260]^x[261]^x[262]^x[264]^x[266]^x[268]^x[269]^x[273]^x[275]^x[276]^x[282]^x[285]^x[286]^x[287]^x[288]^x[289]^x[291]^x[292]^x[293]^x[294]^x[297]^u[61]^u[57]^u[55]^u[53]^u[51]^u[48]^u[46]^u[45]^u[42]^u[41]^u[39]^u[38]^u[37]^u[35]^u[33]^u[31]^u[30]^u[26]^u[24]^u[23]^u[17]^u[14]^u[13]^u[12]^u[11]^u[10]^u[8]^u[7]^u[6]^u[5]^u[2];
	y[117] = x[53]^x[239]^x[243]^x[245]^x[247]^x[249]^x[252]^x[254]^x[255]^x[258]^x[259]^x[261]^x[262]^x[263]^x[265]^x[267]^x[269]^x[270]^x[274]^x[276]^x[277]^x[283]^x[286]^x[287]^x[288]^x[289]^x[290]^x[292]^x[293]^x[294]^x[295]^x[298]^u[60]^u[56]^u[54]^u[52]^u[50]^u[47]^u[45]^u[44]^u[41]^u[40]^u[38]^u[37]^u[36]^u[34]^u[32]^u[30]^u[29]^u[25]^u[23]^u[22]^u[16]^u[13]^u[12]^u[11]^u[10]^u[9]^u[7]^u[6]^u[5]^u[4]^u[1];
	y[118] = x[54]^x[240]^x[244]^x[246]^x[248]^x[250]^x[253]^x[255]^x[256]^x[259]^x[260]^x[262]^x[263]^x[264]^x[266]^x[268]^x[270]^x[271]^x[275]^x[277]^x[278]^x[284]^x[287]^x[288]^x[289]^x[290]^x[291]^x[293]^x[294]^x[295]^x[296]^x[299]^u[59]^u[55]^u[53]^u[51]^u[49]^u[46]^u[44]^u[43]^u[40]^u[39]^u[37]^u[36]^u[35]^u[33]^u[31]^u[29]^u[28]^u[24]^u[22]^u[21]^u[15]^u[12]^u[11]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4]^u[3]^u[0];
	y[119] = x[55]^x[241]^x[245]^x[247]^x[249]^x[251]^x[254]^x[256]^x[257]^x[260]^x[261]^x[263]^x[264]^x[265]^x[267]^x[269]^x[271]^x[272]^x[276]^x[278]^x[279]^x[285]^x[288]^x[289]^x[290]^x[291]^x[292]^x[294]^x[295]^x[296]^x[297]^u[58]^u[54]^u[52]^u[50]^u[48]^u[45]^u[43]^u[42]^u[39]^u[38]^u[36]^u[35]^u[34]^u[32]^u[30]^u[28]^u[27]^u[23]^u[21]^u[20]^u[14]^u[11]^u[10]^u[9]^u[8]^u[7]^u[5]^u[4]^u[3]^u[2];
	y[120] = x[56]^x[236]^x[238]^x[239]^x[241]^x[242]^x[245]^x[246]^x[248]^x[250]^x[252]^x[257]^x[258]^x[260]^x[261]^x[262]^x[265]^x[266]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[276]^x[277]^x[285]^x[286]^x[287]^x[290]^x[291]^x[294]^x[296]^x[297]^u[63]^u[61]^u[60]^u[58]^u[57]^u[54]^u[53]^u[51]^u[49]^u[47]^u[42]^u[41]^u[39]^u[38]^u[37]^u[34]^u[33]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[23]^u[22]^u[14]^u[13]^u[12]^u[9]^u[8]^u[5]^u[3]^u[2];
	y[121] = x[57]^x[236]^x[237]^x[238]^x[240]^x[241]^x[242]^x[243]^x[245]^x[246]^x[247]^x[249]^x[251]^x[253]^x[255]^x[258]^x[259]^x[260]^x[261]^x[262]^x[263]^x[264]^x[266]^x[267]^x[270]^x[272]^x[273]^x[274]^x[276]^x[277]^x[278]^x[279]^x[280]^x[285]^x[286]^x[288]^x[289]^x[291]^x[293]^x[294]^x[297]^u[63]^u[62]^u[61]^u[59]^u[58]^u[57]^u[56]^u[54]^u[53]^u[52]^u[50]^u[48]^u[46]^u[44]^u[41]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[33]^u[32]^u[29]^u[27]^u[26]^u[25]^u[23]^u[22]^u[21]^u[20]^u[19]^u[14]^u[13]^u[11]^u[10]^u[8]^u[6]^u[5]^u[2];
	y[122] = x[58]^x[237]^x[238]^x[239]^x[241]^x[242]^x[243]^x[244]^x[246]^x[247]^x[248]^x[250]^x[252]^x[254]^x[256]^x[259]^x[260]^x[261]^x[262]^x[263]^x[264]^x[265]^x[267]^x[268]^x[271]^x[273]^x[274]^x[275]^x[277]^x[278]^x[279]^x[280]^x[281]^x[286]^x[287]^x[289]^x[290]^x[292]^x[294]^x[295]^x[298]^u[62]^u[61]^u[60]^u[58]^u[57]^u[56]^u[55]^u[53]^u[52]^u[51]^u[49]^u[47]^u[45]^u[43]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[32]^u[31]^u[28]^u[26]^u[25]^u[24]^u[22]^u[21]^u[20]^u[19]^u[18]^u[13]^u[12]^u[10]^u[9]^u[7]^u[5]^u[4]^u[1];
	y[123] = x[59]^x[238]^x[239]^x[240]^x[242]^x[243]^x[244]^x[245]^x[247]^x[248]^x[249]^x[251]^x[253]^x[255]^x[257]^x[260]^x[261]^x[262]^x[263]^x[264]^x[265]^x[266]^x[268]^x[269]^x[272]^x[274]^x[275]^x[276]^x[278]^x[279]^x[280]^x[281]^x[282]^x[287]^x[288]^x[290]^x[291]^x[293]^x[295]^x[296]^x[299]^u[61]^u[60]^u[59]^u[57]^u[56]^u[55]^u[54]^u[52]^u[51]^u[50]^u[48]^u[46]^u[44]^u[42]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[31]^u[30]^u[27]^u[25]^u[24]^u[23]^u[21]^u[20]^u[19]^u[18]^u[17]^u[12]^u[11]^u[9]^u[8]^u[6]^u[4]^u[3]^u[0];
	y[124] = x[60]^x[239]^x[240]^x[241]^x[243]^x[244]^x[245]^x[246]^x[248]^x[249]^x[250]^x[252]^x[254]^x[256]^x[258]^x[261]^x[262]^x[263]^x[264]^x[265]^x[266]^x[267]^x[269]^x[270]^x[273]^x[275]^x[276]^x[277]^x[279]^x[280]^x[281]^x[282]^x[283]^x[288]^x[289]^x[291]^x[292]^x[294]^x[296]^x[297]^u[60]^u[59]^u[58]^u[56]^u[55]^u[54]^u[53]^u[51]^u[50]^u[49]^u[47]^u[45]^u[43]^u[41]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32]^u[30]^u[29]^u[26]^u[24]^u[23]^u[22]^u[20]^u[19]^u[18]^u[17]^u[16]^u[11]^u[10]^u[8]^u[7]^u[5]^u[3]^u[2];
	y[125] = x[61]^x[240]^x[241]^x[242]^x[244]^x[245]^x[246]^x[247]^x[249]^x[250]^x[251]^x[253]^x[255]^x[257]^x[259]^x[262]^x[263]^x[264]^x[265]^x[266]^x[267]^x[268]^x[270]^x[271]^x[274]^x[276]^x[277]^x[278]^x[280]^x[281]^x[282]^x[283]^x[284]^x[289]^x[290]^x[292]^x[293]^x[295]^x[297]^x[298]^u[59]^u[58]^u[57]^u[55]^u[54]^u[53]^u[52]^u[50]^u[49]^u[48]^u[46]^u[44]^u[42]^u[40]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32]^u[31]^u[29]^u[28]^u[25]^u[23]^u[22]^u[21]^u[19]^u[18]^u[17]^u[16]^u[15]^u[10]^u[9]^u[7]^u[6]^u[4]^u[2]^u[1];
	y[126] = x[62]^x[236]^x[238]^x[239]^x[242]^x[243]^x[246]^x[247]^x[248]^x[250]^x[251]^x[252]^x[254]^x[255]^x[256]^x[258]^x[263]^x[265]^x[266]^x[267]^x[268]^x[272]^x[275]^x[276]^x[277]^x[278]^x[280]^x[281]^x[282]^x[283]^x[284]^x[287]^x[289]^x[290]^x[291]^x[292]^x[295]^x[296]^x[299]^u[63]^u[61]^u[60]^u[57]^u[56]^u[53]^u[52]^u[51]^u[49]^u[48]^u[47]^u[45]^u[44]^u[43]^u[41]^u[36]^u[34]^u[33]^u[32]^u[31]^u[27]^u[24]^u[23]^u[22]^u[21]^u[19]^u[18]^u[17]^u[16]^u[15]^u[12]^u[10]^u[9]^u[8]^u[7]^u[4]^u[3]^u[0];
	y[127] = x[63]^x[237]^x[239]^x[240]^x[243]^x[244]^x[247]^x[248]^x[249]^x[251]^x[252]^x[253]^x[255]^x[256]^x[257]^x[259]^x[264]^x[266]^x[267]^x[268]^x[269]^x[273]^x[276]^x[277]^x[278]^x[279]^x[281]^x[282]^x[283]^x[284]^x[285]^x[288]^x[290]^x[291]^x[292]^x[293]^x[296]^x[297]^u[62]^u[60]^u[59]^u[56]^u[55]^u[52]^u[51]^u[50]^u[48]^u[47]^u[46]^u[44]^u[43]^u[42]^u[40]^u[35]^u[33]^u[32]^u[31]^u[30]^u[26]^u[23]^u[22]^u[21]^u[20]^u[18]^u[17]^u[16]^u[15]^u[14]^u[11]^u[9]^u[8]^u[7]^u[6]^u[3]^u[2];
	y[128] = x[64]^x[236]^x[239]^x[240]^x[244]^x[248]^x[249]^x[250]^x[252]^x[253]^x[254]^x[255]^x[256]^x[257]^x[258]^x[264]^x[265]^x[267]^x[268]^x[270]^x[271]^x[274]^x[276]^x[277]^x[278]^x[282]^x[283]^x[284]^x[286]^x[287]^x[291]^x[295]^x[297]^u[63]^u[60]^u[59]^u[55]^u[51]^u[50]^u[49]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[35]^u[34]^u[32]^u[31]^u[29]^u[28]^u[25]^u[23]^u[22]^u[21]^u[17]^u[16]^u[15]^u[13]^u[12]^u[8]^u[4]^u[2];
	y[129] = x[65]^x[237]^x[240]^x[241]^x[245]^x[249]^x[250]^x[251]^x[253]^x[254]^x[255]^x[256]^x[257]^x[258]^x[259]^x[265]^x[266]^x[268]^x[269]^x[271]^x[272]^x[275]^x[277]^x[278]^x[279]^x[283]^x[284]^x[285]^x[287]^x[288]^x[292]^x[296]^x[298]^u[62]^u[59]^u[58]^u[54]^u[50]^u[49]^u[48]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40]^u[34]^u[33]^u[31]^u[30]^u[28]^u[27]^u[24]^u[22]^u[21]^u[20]^u[16]^u[15]^u[14]^u[12]^u[11]^u[7]^u[3]^u[1];
	y[130] = x[66]^x[238]^x[241]^x[242]^x[246]^x[250]^x[251]^x[252]^x[254]^x[255]^x[256]^x[257]^x[258]^x[259]^x[260]^x[266]^x[267]^x[269]^x[270]^x[272]^x[273]^x[276]^x[278]^x[279]^x[280]^x[284]^x[285]^x[286]^x[288]^x[289]^x[293]^x[297]^x[299]^u[61]^u[58]^u[57]^u[53]^u[49]^u[48]^u[47]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40]^u[39]^u[33]^u[32]^u[30]^u[29]^u[27]^u[26]^u[23]^u[21]^u[20]^u[19]^u[15]^u[14]^u[13]^u[11]^u[10]^u[6]^u[2]^u[0];
	y[131] = x[67]^x[236]^x[238]^x[241]^x[242]^x[243]^x[245]^x[247]^x[251]^x[252]^x[253]^x[256]^x[257]^x[258]^x[259]^x[261]^x[264]^x[267]^x[268]^x[269]^x[270]^x[273]^x[274]^x[276]^x[277]^x[281]^x[286]^x[290]^x[292]^x[293]^x[295]^u[63]^u[61]^u[58]^u[57]^u[56]^u[54]^u[52]^u[48]^u[47]^u[46]^u[43]^u[42]^u[41]^u[40]^u[38]^u[35]^u[32]^u[31]^u[30]^u[29]^u[26]^u[25]^u[23]^u[22]^u[18]^u[13]^u[9]^u[7]^u[6]^u[4];
	y[132] = x[68]^x[236]^x[237]^x[238]^x[241]^x[242]^x[243]^x[244]^x[245]^x[246]^x[248]^x[252]^x[253]^x[254]^x[255]^x[257]^x[258]^x[259]^x[262]^x[264]^x[265]^x[268]^x[270]^x[274]^x[275]^x[276]^x[277]^x[278]^x[279]^x[280]^x[282]^x[285]^x[289]^x[291]^x[292]^x[295]^x[296]^x[298]^u[63]^u[62]^u[61]^u[58]^u[57]^u[56]^u[55]^u[54]^u[53]^u[51]^u[47]^u[46]^u[45]^u[44]^u[42]^u[41]^u[40]^u[37]^u[35]^u[34]^u[31]^u[29]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[17]^u[14]^u[10]^u[8]^u[7]^u[4]^u[3]^u[1];
	y[133] = x[69]^x[237]^x[238]^x[239]^x[242]^x[243]^x[244]^x[245]^x[246]^x[247]^x[249]^x[253]^x[254]^x[255]^x[256]^x[258]^x[259]^x[260]^x[263]^x[265]^x[266]^x[269]^x[271]^x[275]^x[276]^x[277]^x[278]^x[279]^x[280]^x[281]^x[283]^x[286]^x[290]^x[292]^x[293]^x[296]^x[297]^x[299]^u[62]^u[61]^u[60]^u[57]^u[56]^u[55]^u[54]^u[53]^u[52]^u[50]^u[46]^u[45]^u[44]^u[43]^u[41]^u[40]^u[39]^u[36]^u[34]^u[33]^u[30]^u[28]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[16]^u[13]^u[9]^u[7]^u[6]^u[3]^u[2]^u[0];
	y[134] = x[70]^x[236]^x[240]^x[241]^x[243]^x[244]^x[246]^x[247]^x[248]^x[250]^x[254]^x[256]^x[257]^x[259]^x[261]^x[266]^x[267]^x[269]^x[270]^x[271]^x[272]^x[277]^x[278]^x[281]^x[282]^x[284]^x[285]^x[289]^x[291]^x[292]^x[295]^x[297]^u[63]^u[59]^u[58]^u[56]^u[55]^u[53]^u[52]^u[51]^u[49]^u[45]^u[43]^u[42]^u[40]^u[38]^u[33]^u[32]^u[30]^u[29]^u[28]^u[27]^u[22]^u[21]^u[18]^u[17]^u[15]^u[14]^u[10]^u[8]^u[7]^u[4]^u[2];
	y[135] = x[71]^x[236]^x[237]^x[238]^x[239]^x[242]^x[244]^x[247]^x[248]^x[249]^x[251]^x[257]^x[258]^x[262]^x[264]^x[267]^x[268]^x[269]^x[270]^x[272]^x[273]^x[276]^x[278]^x[280]^x[282]^x[283]^x[286]^x[287]^x[289]^x[290]^x[294]^x[295]^x[296]^u[63]^u[62]^u[61]^u[60]^u[57]^u[55]^u[52]^u[51]^u[50]^u[48]^u[42]^u[41]^u[37]^u[35]^u[32]^u[31]^u[30]^u[29]^u[27]^u[26]^u[23]^u[21]^u[19]^u[17]^u[16]^u[13]^u[12]^u[10]^u[9]^u[5]^u[4]^u[3];
	y[136] = x[72]^x[237]^x[238]^x[239]^x[240]^x[243]^x[245]^x[248]^x[249]^x[250]^x[252]^x[258]^x[259]^x[263]^x[265]^x[268]^x[269]^x[270]^x[271]^x[273]^x[274]^x[277]^x[279]^x[281]^x[283]^x[284]^x[287]^x[288]^x[290]^x[291]^x[295]^x[296]^x[297]^u[62]^u[61]^u[60]^u[59]^u[56]^u[54]^u[51]^u[50]^u[49]^u[47]^u[41]^u[40]^u[36]^u[34]^u[31]^u[30]^u[29]^u[28]^u[26]^u[25]^u[22]^u[20]^u[18]^u[16]^u[15]^u[12]^u[11]^u[9]^u[8]^u[4]^u[3]^u[2];
	y[137] = x[73]^x[236]^x[240]^x[244]^x[245]^x[246]^x[249]^x[250]^x[251]^x[253]^x[255]^x[259]^x[266]^x[270]^x[272]^x[274]^x[275]^x[276]^x[278]^x[279]^x[282]^x[284]^x[287]^x[288]^x[291]^x[293]^x[294]^x[295]^x[296]^x[297]^u[63]^u[59]^u[55]^u[54]^u[53]^u[50]^u[49]^u[48]^u[46]^u[44]^u[40]^u[33]^u[29]^u[27]^u[25]^u[24]^u[23]^u[21]^u[20]^u[17]^u[15]^u[12]^u[11]^u[8]^u[6]^u[5]^u[4]^u[3]^u[2];
	y[138] = x[74]^x[237]^x[241]^x[245]^x[246]^x[247]^x[250]^x[251]^x[252]^x[254]^x[256]^x[260]^x[267]^x[271]^x[273]^x[275]^x[276]^x[277]^x[279]^x[280]^x[283]^x[285]^x[288]^x[289]^x[292]^x[294]^x[295]^x[296]^x[297]^x[298]^u[62]^u[58]^u[54]^u[53]^u[52]^u[49]^u[48]^u[47]^u[45]^u[43]^u[39]^u[32]^u[28]^u[26]^u[24]^u[23]^u[22]^u[20]^u[19]^u[16]^u[14]^u[11]^u[10]^u[7]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[139] = x[75]^x[238]^x[242]^x[246]^x[247]^x[248]^x[251]^x[252]^x[253]^x[255]^x[257]^x[261]^x[268]^x[272]^x[274]^x[276]^x[277]^x[278]^x[280]^x[281]^x[284]^x[286]^x[289]^x[290]^x[293]^x[295]^x[296]^x[297]^x[298]^x[299]^u[61]^u[57]^u[53]^u[52]^u[51]^u[48]^u[47]^u[46]^u[44]^u[42]^u[38]^u[31]^u[27]^u[25]^u[23]^u[22]^u[21]^u[19]^u[18]^u[15]^u[13]^u[10]^u[9]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[140] = x[76]^x[236]^x[238]^x[241]^x[243]^x[245]^x[247]^x[248]^x[249]^x[252]^x[253]^x[254]^x[255]^x[256]^x[258]^x[260]^x[262]^x[264]^x[271]^x[273]^x[275]^x[276]^x[277]^x[278]^x[280]^x[281]^x[282]^x[289]^x[290]^x[291]^x[292]^x[293]^x[295]^x[296]^x[297]^x[299]^u[63]^u[61]^u[58]^u[56]^u[54]^u[52]^u[51]^u[50]^u[47]^u[46]^u[45]^u[44]^u[43]^u[41]^u[39]^u[37]^u[35]^u[28]^u[26]^u[24]^u[23]^u[22]^u[21]^u[19]^u[18]^u[17]^u[10]^u[9]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[0];
	y[141] = x[77]^x[236]^x[237]^x[238]^x[241]^x[242]^x[244]^x[245]^x[246]^x[248]^x[249]^x[250]^x[253]^x[254]^x[256]^x[257]^x[259]^x[260]^x[261]^x[263]^x[264]^x[265]^x[269]^x[271]^x[272]^x[274]^x[277]^x[278]^x[280]^x[281]^x[282]^x[283]^x[285]^x[287]^x[289]^x[290]^x[291]^x[295]^x[296]^x[297]^u[63]^u[62]^u[61]^u[58]^u[57]^u[55]^u[54]^u[53]^u[51]^u[50]^u[49]^u[46]^u[45]^u[43]^u[42]^u[40]^u[39]^u[38]^u[36]^u[35]^u[34]^u[30]^u[28]^u[27]^u[25]^u[22]^u[21]^u[19]^u[18]^u[17]^u[16]^u[14]^u[12]^u[10]^u[9]^u[8]^u[4]^u[3]^u[2];
	y[142] = x[78]^x[237]^x[238]^x[239]^x[242]^x[243]^x[245]^x[246]^x[247]^x[249]^x[250]^x[251]^x[254]^x[255]^x[257]^x[258]^x[260]^x[261]^x[262]^x[264]^x[265]^x[266]^x[270]^x[272]^x[273]^x[275]^x[278]^x[279]^x[281]^x[282]^x[283]^x[284]^x[286]^x[288]^x[290]^x[291]^x[292]^x[296]^x[297]^x[298]^u[62]^u[61]^u[60]^u[57]^u[56]^u[54]^u[53]^u[52]^u[50]^u[49]^u[48]^u[45]^u[44]^u[42]^u[41]^u[39]^u[38]^u[37]^u[35]^u[34]^u[33]^u[29]^u[27]^u[26]^u[24]^u[21]^u[20]^u[18]^u[17]^u[16]^u[15]^u[13]^u[11]^u[9]^u[8]^u[7]^u[3]^u[2]^u[1];
	y[143] = x[79]^x[236]^x[240]^x[241]^x[243]^x[244]^x[245]^x[246]^x[247]^x[248]^x[250]^x[251]^x[252]^x[256]^x[258]^x[259]^x[260]^x[261]^x[262]^x[263]^x[264]^x[265]^x[266]^x[267]^x[269]^x[273]^x[274]^x[282]^x[283]^x[284]^x[291]^x[294]^x[295]^x[297]^x[299]^u[63]^u[59]^u[58]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[49]^u[48]^u[47]^u[43]^u[41]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32]^u[30]^u[26]^u[25]^u[17]^u[16]^u[15]^u[8]^u[5]^u[4]^u[2]^u[0];
	y[144] = x[80]^x[236]^x[237]^x[238]^x[239]^x[242]^x[244]^x[246]^x[247]^x[248]^x[249]^x[251]^x[252]^x[253]^x[255]^x[257]^x[259]^x[261]^x[262]^x[263]^x[265]^x[266]^x[267]^x[268]^x[269]^x[270]^x[271]^x[274]^x[275]^x[276]^x[279]^x[280]^x[283]^x[284]^x[287]^x[289]^x[293]^x[294]^x[296]^u[63]^u[62]^u[61]^u[60]^u[57]^u[55]^u[53]^u[52]^u[51]^u[50]^u[48]^u[47]^u[46]^u[44]^u[42]^u[40]^u[38]^u[37]^u[36]^u[34]^u[33]^u[32]^u[31]^u[30]^u[29]^u[28]^u[25]^u[24]^u[23]^u[20]^u[19]^u[16]^u[15]^u[12]^u[10]^u[6]^u[5]^u[3];
	y[145] = x[81]^x[237]^x[238]^x[239]^x[240]^x[243]^x[245]^x[247]^x[248]^x[249]^x[250]^x[252]^x[253]^x[254]^x[256]^x[258]^x[260]^x[262]^x[263]^x[264]^x[266]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[275]^x[276]^x[277]^x[280]^x[281]^x[284]^x[285]^x[288]^x[290]^x[294]^x[295]^x[297]^u[62]^u[61]^u[60]^u[59]^u[56]^u[54]^u[52]^u[51]^u[50]^u[49]^u[47]^u[46]^u[45]^u[43]^u[41]^u[39]^u[37]^u[36]^u[35]^u[33]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[24]^u[23]^u[22]^u[19]^u[18]^u[15]^u[14]^u[11]^u[9]^u[5]^u[4]^u[2];
	y[146] = x[82]^x[238]^x[239]^x[240]^x[241]^x[244]^x[246]^x[248]^x[249]^x[250]^x[251]^x[253]^x[254]^x[255]^x[257]^x[259]^x[261]^x[263]^x[264]^x[265]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[276]^x[277]^x[278]^x[281]^x[282]^x[285]^x[286]^x[289]^x[291]^x[295]^x[296]^x[298]^u[61]^u[60]^u[59]^u[58]^u[55]^u[53]^u[51]^u[50]^u[49]^u[48]^u[46]^u[45]^u[44]^u[42]^u[40]^u[38]^u[36]^u[35]^u[34]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[23]^u[22]^u[21]^u[18]^u[17]^u[14]^u[13]^u[10]^u[8]^u[4]^u[3]^u[1];
	y[147] = x[83]^x[236]^x[238]^x[240]^x[242]^x[247]^x[249]^x[250]^x[251]^x[252]^x[254]^x[256]^x[258]^x[262]^x[265]^x[266]^x[268]^x[270]^x[272]^x[273]^x[274]^x[276]^x[277]^x[278]^x[280]^x[282]^x[283]^x[285]^x[286]^x[289]^x[290]^x[293]^x[294]^x[295]^x[296]^x[297]^x[298]^x[299]^u[63]^u[61]^u[59]^u[57]^u[52]^u[50]^u[49]^u[48]^u[47]^u[45]^u[43]^u[41]^u[37]^u[34]^u[33]^u[31]^u[29]^u[27]^u[26]^u[25]^u[23]^u[22]^u[21]^u[19]^u[17]^u[16]^u[14]^u[13]^u[10]^u[9]^u[6]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[148] = x[84]^x[236]^x[237]^x[238]^x[243]^x[245]^x[248]^x[250]^x[251]^x[252]^x[253]^x[257]^x[259]^x[260]^x[263]^x[264]^x[266]^x[267]^x[273]^x[274]^x[275]^x[276]^x[277]^x[278]^x[280]^x[281]^x[283]^x[284]^x[285]^x[286]^x[289]^x[290]^x[291]^x[292]^x[293]^x[296]^x[297]^x[299]^u[63]^u[62]^u[61]^u[56]^u[54]^u[51]^u[49]^u[48]^u[47]^u[46]^u[42]^u[40]^u[39]^u[36]^u[35]^u[33]^u[32]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[19]^u[18]^u[16]^u[15]^u[14]^u[13]^u[10]^u[9]^u[8]^u[7]^u[6]^u[3]^u[2]^u[0];
	y[149] = x[85]^x[236]^x[237]^x[241]^x[244]^x[245]^x[246]^x[249]^x[251]^x[252]^x[253]^x[254]^x[255]^x[258]^x[261]^x[265]^x[267]^x[268]^x[269]^x[271]^x[274]^x[275]^x[277]^x[278]^x[280]^x[281]^x[282]^x[284]^x[286]^x[289]^x[290]^x[291]^x[295]^x[297]^u[63]^u[62]^u[58]^u[55]^u[54]^u[53]^u[50]^u[48]^u[47]^u[46]^u[45]^u[44]^u[41]^u[38]^u[34]^u[32]^u[31]^u[30]^u[28]^u[25]^u[24]^u[22]^u[21]^u[19]^u[18]^u[17]^u[15]^u[13]^u[10]^u[9]^u[8]^u[4]^u[2];
	y[150] = x[86]^x[236]^x[237]^x[239]^x[241]^x[242]^x[246]^x[247]^x[250]^x[252]^x[253]^x[254]^x[256]^x[259]^x[260]^x[262]^x[264]^x[266]^x[268]^x[270]^x[271]^x[272]^x[275]^x[278]^x[280]^x[281]^x[282]^x[283]^x[289]^x[290]^x[291]^x[293]^x[294]^x[295]^x[296]^u[63]^u[62]^u[60]^u[58]^u[57]^u[53]^u[52]^u[49]^u[47]^u[46]^u[45]^u[43]^u[40]^u[39]^u[37]^u[35]^u[33]^u[31]^u[29]^u[28]^u[27]^u[24]^u[21]^u[19]^u[18]^u[17]^u[16]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4]^u[3];
	y[151] = x[87]^x[237]^x[238]^x[240]^x[242]^x[243]^x[247]^x[248]^x[251]^x[253]^x[254]^x[255]^x[257]^x[260]^x[261]^x[263]^x[265]^x[267]^x[269]^x[271]^x[272]^x[273]^x[276]^x[279]^x[281]^x[282]^x[283]^x[284]^x[290]^x[291]^x[292]^x[294]^x[295]^x[296]^x[297]^u[62]^u[61]^u[59]^u[57]^u[56]^u[52]^u[51]^u[48]^u[46]^u[45]^u[44]^u[42]^u[39]^u[38]^u[36]^u[34]^u[32]^u[30]^u[28]^u[27]^u[26]^u[23]^u[20]^u[18]^u[17]^u[16]^u[15]^u[9]^u[8]^u[7]^u[5]^u[4]^u[3]^u[2];
	y[152] = x[88]^x[238]^x[239]^x[241]^x[243]^x[244]^x[248]^x[249]^x[252]^x[254]^x[255]^x[256]^x[258]^x[261]^x[262]^x[264]^x[266]^x[268]^x[270]^x[272]^x[273]^x[274]^x[277]^x[280]^x[282]^x[283]^x[284]^x[285]^x[291]^x[292]^x[293]^x[295]^x[296]^x[297]^x[298]^u[61]^u[60]^u[58]^u[56]^u[55]^u[51]^u[50]^u[47]^u[45]^u[44]^u[43]^u[41]^u[38]^u[37]^u[35]^u[33]^u[31]^u[29]^u[27]^u[26]^u[25]^u[22]^u[19]^u[17]^u[16]^u[15]^u[14]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1];
	y[153] = x[89]^x[236]^x[238]^x[240]^x[241]^x[242]^x[244]^x[249]^x[250]^x[253]^x[256]^x[257]^x[259]^x[260]^x[262]^x[263]^x[264]^x[265]^x[267]^x[273]^x[274]^x[275]^x[276]^x[278]^x[279]^x[280]^x[281]^x[283]^x[284]^x[286]^x[287]^x[289]^x[295]^x[296]^x[297]^x[299]^u[63]^u[61]^u[59]^u[58]^u[57]^u[55]^u[50]^u[49]^u[46]^u[43]^u[42]^u[40]^u[39]^u[37]^u[36]^u[35]^u[34]^u[32]^u[26]^u[25]^u[24]^u[23]^u[21]^u[20]^u[19]^u[18]^u[16]^u[15]^u[13]^u[12]^u[10]^u[4]^u[3]^u[2]^u[0];
	y[154] = x[90]^x[236]^x[237]^x[238]^x[242]^x[243]^x[250]^x[251]^x[254]^x[255]^x[257]^x[258]^x[261]^x[263]^x[265]^x[266]^x[268]^x[269]^x[271]^x[274]^x[275]^x[277]^x[281]^x[282]^x[284]^x[288]^x[289]^x[290]^x[292]^x[293]^x[294]^x[295]^x[296]^x[297]^u[63]^u[62]^u[61]^u[57]^u[56]^u[49]^u[48]^u[45]^u[44]^u[42]^u[41]^u[38]^u[36]^u[34]^u[33]^u[31]^u[30]^u[28]^u[25]^u[24]^u[22]^u[18]^u[17]^u[15]^u[11]^u[10]^u[9]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2];
	y[155] = x[91]^x[236]^x[237]^x[241]^x[243]^x[244]^x[245]^x[251]^x[252]^x[256]^x[258]^x[259]^x[260]^x[262]^x[266]^x[267]^x[270]^x[271]^x[272]^x[275]^x[278]^x[279]^x[280]^x[282]^x[283]^x[287]^x[290]^x[291]^x[292]^x[296]^x[297]^u[63]^u[62]^u[58]^u[56]^u[55]^u[54]^u[48]^u[47]^u[43]^u[41]^u[40]^u[39]^u[37]^u[33]^u[32]^u[29]^u[28]^u[27]^u[24]^u[21]^u[20]^u[19]^u[17]^u[16]^u[12]^u[9]^u[8]^u[7]^u[3]^u[2];
	y[156] = x[92]^x[236]^x[237]^x[239]^x[241]^x[242]^x[244]^x[246]^x[252]^x[253]^x[255]^x[257]^x[259]^x[261]^x[263]^x[264]^x[267]^x[268]^x[269]^x[272]^x[273]^x[281]^x[283]^x[284]^x[285]^x[287]^x[288]^x[289]^x[291]^x[294]^x[295]^x[297]^u[63]^u[62]^u[60]^u[58]^u[57]^u[55]^u[53]^u[47]^u[46]^u[44]^u[42]^u[40]^u[38]^u[36]^u[35]^u[32]^u[31]^u[30]^u[27]^u[26]^u[18]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[8]^u[5]^u[4]^u[2];
	y[157] = x[93]^x[237]^x[238]^x[240]^x[242]^x[243]^x[245]^x[247]^x[253]^x[254]^x[256]^x[258]^x[260]^x[262]^x[264]^x[265]^x[268]^x[269]^x[270]^x[273]^x[274]^x[282]^x[284]^x[285]^x[286]^x[288]^x[289]^x[290]^x[292]^x[295]^x[296]^x[298]^u[62]^u[61]^u[59]^u[57]^u[56]^u[54]^u[52]^u[46]^u[45]^u[43]^u[41]^u[39]^u[37]^u[35]^u[34]^u[31]^u[30]^u[29]^u[26]^u[25]^u[17]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[7]^u[4]^u[3]^u[1];
	y[158] = x[94]^x[238]^x[239]^x[241]^x[243]^x[244]^x[246]^x[248]^x[254]^x[255]^x[257]^x[259]^x[261]^x[263]^x[265]^x[266]^x[269]^x[270]^x[271]^x[274]^x[275]^x[283]^x[285]^x[286]^x[287]^x[289]^x[290]^x[291]^x[293]^x[296]^x[297]^x[299]^u[61]^u[60]^u[58]^u[56]^u[55]^u[53]^u[51]^u[45]^u[44]^u[42]^u[40]^u[38]^u[36]^u[34]^u[33]^u[30]^u[29]^u[28]^u[25]^u[24]^u[16]^u[14]^u[13]^u[12]^u[10]^u[9]^u[8]^u[6]^u[3]^u[2]^u[0];
	y[159] = x[95]^x[236]^x[238]^x[240]^x[241]^x[242]^x[244]^x[247]^x[249]^x[256]^x[258]^x[262]^x[266]^x[267]^x[269]^x[270]^x[272]^x[275]^x[279]^x[280]^x[284]^x[285]^x[286]^x[288]^x[289]^x[290]^x[291]^x[293]^x[295]^x[297]^u[63]^u[61]^u[59]^u[58]^u[57]^u[55]^u[52]^u[50]^u[43]^u[41]^u[37]^u[33]^u[32]^u[30]^u[29]^u[27]^u[24]^u[20]^u[19]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[6]^u[4]^u[2];
	y[160] = x[96]^x[237]^x[239]^x[241]^x[242]^x[243]^x[245]^x[248]^x[250]^x[257]^x[259]^x[263]^x[267]^x[268]^x[270]^x[271]^x[273]^x[276]^x[280]^x[281]^x[285]^x[286]^x[287]^x[289]^x[290]^x[291]^x[292]^x[294]^x[296]^x[298]^u[62]^u[60]^u[58]^u[57]^u[56]^u[54]^u[51]^u[49]^u[42]^u[40]^u[36]^u[32]^u[31]^u[29]^u[28]^u[26]^u[23]^u[19]^u[18]^u[14]^u[13]^u[12]^u[10]^u[9]^u[8]^u[7]^u[5]^u[3]^u[1];
	y[161] = x[97]^x[238]^x[240]^x[242]^x[243]^x[244]^x[246]^x[249]^x[251]^x[258]^x[260]^x[264]^x[268]^x[269]^x[271]^x[272]^x[274]^x[277]^x[281]^x[282]^x[286]^x[287]^x[288]^x[290]^x[291]^x[292]^x[293]^x[295]^x[297]^x[299]^u[61]^u[59]^u[57]^u[56]^u[55]^u[53]^u[50]^u[48]^u[41]^u[39]^u[35]^u[31]^u[30]^u[28]^u[27]^u[25]^u[22]^u[18]^u[17]^u[13]^u[12]^u[11]^u[9]^u[8]^u[7]^u[6]^u[4]^u[2]^u[0];
	y[162] = x[98]^x[239]^x[241]^x[243]^x[244]^x[245]^x[247]^x[250]^x[252]^x[259]^x[261]^x[265]^x[269]^x[270]^x[272]^x[273]^x[275]^x[278]^x[282]^x[283]^x[287]^x[288]^x[289]^x[291]^x[292]^x[293]^x[294]^x[296]^x[298]^u[60]^u[58]^u[56]^u[55]^u[54]^u[52]^u[49]^u[47]^u[40]^u[38]^u[34]^u[30]^u[29]^u[27]^u[26]^u[24]^u[21]^u[17]^u[16]^u[12]^u[11]^u[10]^u[8]^u[7]^u[6]^u[5]^u[3]^u[1];
	y[163] = x[99]^x[240]^x[242]^x[244]^x[245]^x[246]^x[248]^x[251]^x[253]^x[260]^x[262]^x[266]^x[270]^x[271]^x[273]^x[274]^x[276]^x[279]^x[283]^x[284]^x[288]^x[289]^x[290]^x[292]^x[293]^x[294]^x[295]^x[297]^x[299]^u[59]^u[57]^u[55]^u[54]^u[53]^u[51]^u[48]^u[46]^u[39]^u[37]^u[33]^u[29]^u[28]^u[26]^u[25]^u[23]^u[20]^u[16]^u[15]^u[11]^u[10]^u[9]^u[7]^u[6]^u[5]^u[4]^u[2]^u[0];
	y[164] = x[100]^x[241]^x[243]^x[245]^x[246]^x[247]^x[249]^x[252]^x[254]^x[261]^x[263]^x[267]^x[271]^x[272]^x[274]^x[275]^x[277]^x[280]^x[284]^x[285]^x[289]^x[290]^x[291]^x[293]^x[294]^x[295]^x[296]^x[298]^u[58]^u[56]^u[54]^u[53]^u[52]^u[50]^u[47]^u[45]^u[38]^u[36]^u[32]^u[28]^u[27]^u[25]^u[24]^u[22]^u[19]^u[15]^u[14]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4]^u[3]^u[1];
	y[165] = x[101]^x[236]^x[238]^x[239]^x[241]^x[242]^x[244]^x[245]^x[246]^x[247]^x[248]^x[250]^x[253]^x[260]^x[262]^x[268]^x[269]^x[271]^x[272]^x[273]^x[275]^x[278]^x[279]^x[280]^x[281]^x[286]^x[287]^x[289]^x[290]^x[291]^x[293]^x[296]^x[297]^x[298]^x[299]^u[63]^u[61]^u[60]^u[58]^u[57]^u[55]^u[54]^u[53]^u[52]^u[51]^u[49]^u[46]^u[39]^u[37]^u[31]^u[30]^u[28]^u[27]^u[26]^u[24]^u[21]^u[20]^u[19]^u[18]^u[13]^u[12]^u[10]^u[9]^u[8]^u[6]^u[3]^u[2]^u[1]^u[0];
	y[166] = x[102]^x[236]^x[237]^x[238]^x[240]^x[241]^x[242]^x[243]^x[246]^x[247]^x[248]^x[249]^x[251]^x[254]^x[255]^x[260]^x[261]^x[263]^x[264]^x[270]^x[271]^x[272]^x[273]^x[274]^x[281]^x[282]^x[285]^x[288]^x[289]^x[290]^x[291]^x[293]^x[295]^x[297]^x[299]^u[63]^u[62]^u[61]^u[59]^u[58]^u[57]^u[56]^u[53]^u[52]^u[51]^u[50]^u[48]^u[45]^u[44]^u[39]^u[38]^u[36]^u[35]^u[29]^u[28]^u[27]^u[26]^u[25]^u[18]^u[17]^u[14]^u[11]^u[10]^u[9]^u[8]^u[6]^u[4]^u[2]^u[0];
	y[167] = x[103]^x[236]^x[237]^x[242]^x[243]^x[244]^x[245]^x[247]^x[248]^x[249]^x[250]^x[252]^x[256]^x[260]^x[261]^x[262]^x[265]^x[269]^x[272]^x[273]^x[274]^x[275]^x[276]^x[279]^x[280]^x[282]^x[283]^x[285]^x[286]^x[287]^x[290]^x[291]^x[293]^x[295]^x[296]^u[63]^u[62]^u[57]^u[56]^u[55]^u[54]^u[52]^u[51]^u[50]^u[49]^u[47]^u[43]^u[39]^u[38]^u[37]^u[34]^u[30]^u[27]^u[26]^u[25]^u[24]^u[23]^u[20]^u[19]^u[17]^u[16]^u[14]^u[13]^u[12]^u[9]^u[8]^u[6]^u[4]^u[3];
	y[168] = x[104]^x[236]^x[237]^x[239]^x[241]^x[243]^x[244]^x[246]^x[248]^x[249]^x[250]^x[251]^x[253]^x[255]^x[257]^x[260]^x[261]^x[262]^x[263]^x[264]^x[266]^x[269]^x[270]^x[271]^x[273]^x[274]^x[275]^x[277]^x[279]^x[281]^x[283]^x[284]^x[285]^x[286]^x[288]^x[289]^x[291]^x[293]^x[295]^x[296]^x[297]^x[298]^u[63]^u[62]^u[60]^u[58]^u[56]^u[55]^u[53]^u[51]^u[50]^u[49]^u[48]^u[46]^u[44]^u[42]^u[39]^u[38]^u[37]^u[36]^u[35]^u[33]^u[30]^u[29]^u[28]^u[26]^u[25]^u[24]^u[22]^u[20]^u[18]^u[16]^u[15]^u[14]^u[13]^u[11]^u[10]^u[8]^u[6]^u[4]^u[3]^u[2]^u[1];
	y[169] = x[105]^x[236]^x[237]^x[239]^x[240]^x[241]^x[242]^x[244]^x[247]^x[249]^x[250]^x[251]^x[252]^x[254]^x[255]^x[256]^x[258]^x[260]^x[261]^x[262]^x[263]^x[265]^x[267]^x[269]^x[270]^x[272]^x[274]^x[275]^x[278]^x[279]^x[282]^x[284]^x[286]^x[290]^x[293]^x[295]^x[296]^x[297]^x[299]^u[63]^u[62]^u[60]^u[59]^u[58]^u[57]^u[55]^u[52]^u[50]^u[49]^u[48]^u[47]^u[45]^u[44]^u[43]^u[41]^u[39]^u[38]^u[37]^u[36]^u[34]^u[32]^u[30]^u[29]^u[27]^u[25]^u[24]^u[21]^u[20]^u[17]^u[15]^u[13]^u[9]^u[6]^u[4]^u[3]^u[2]^u[0];
	y[170] = x[106]^x[237]^x[238]^x[240]^x[241]^x[242]^x[243]^x[245]^x[248]^x[250]^x[251]^x[252]^x[253]^x[255]^x[256]^x[257]^x[259]^x[261]^x[262]^x[263]^x[264]^x[266]^x[268]^x[270]^x[271]^x[273]^x[275]^x[276]^x[279]^x[280]^x[283]^x[285]^x[287]^x[291]^x[294]^x[296]^x[297]^x[298]^u[62]^u[61]^u[59]^u[58]^u[57]^u[56]^u[54]^u[51]^u[49]^u[48]^u[47]^u[46]^u[44]^u[43]^u[42]^u[40]^u[38]^u[37]^u[36]^u[35]^u[33]^u[31]^u[29]^u[28]^u[26]^u[24]^u[23]^u[20]^u[19]^u[16]^u[14]^u[12]^u[8]^u[5]^u[3]^u[2]^u[1];
	y[171] = x[107]^x[236]^x[242]^x[243]^x[244]^x[245]^x[246]^x[249]^x[251]^x[252]^x[253]^x[254]^x[255]^x[256]^x[257]^x[258]^x[262]^x[263]^x[265]^x[267]^x[272]^x[274]^x[277]^x[279]^x[281]^x[284]^x[285]^x[286]^x[287]^x[288]^x[289]^x[293]^x[294]^x[297]^x[299]^u[63]^u[57]^u[56]^u[55]^u[54]^u[53]^u[50]^u[48]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[37]^u[36]^u[34]^u[32]^u[27]^u[25]^u[22]^u[20]^u[18]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[6]^u[5]^u[2]^u[0];
	y[172] = x[108]^x[237]^x[243]^x[244]^x[245]^x[246]^x[247]^x[250]^x[252]^x[253]^x[254]^x[255]^x[256]^x[257]^x[258]^x[259]^x[263]^x[264]^x[266]^x[268]^x[273]^x[275]^x[278]^x[280]^x[282]^x[285]^x[286]^x[287]^x[288]^x[289]^x[290]^x[294]^x[295]^x[298]^u[62]^u[56]^u[55]^u[54]^u[53]^u[52]^u[49]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40]^u[36]^u[35]^u[33]^u[31]^u[26]^u[24]^u[21]^u[19]^u[17]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[5]^u[4]^u[1];
	y[173] = x[109]^x[236]^x[239]^x[241]^x[244]^x[246]^x[247]^x[248]^x[251]^x[253]^x[254]^x[256]^x[257]^x[258]^x[259]^x[265]^x[267]^x[271]^x[274]^x[280]^x[281]^x[283]^x[285]^x[286]^x[288]^x[290]^x[291]^x[292]^x[293]^x[294]^x[296]^x[298]^x[299]^u[63]^u[60]^u[58]^u[55]^u[53]^u[52]^u[51]^u[48]^u[46]^u[45]^u[43]^u[42]^u[41]^u[40]^u[34]^u[32]^u[28]^u[25]^u[19]^u[18]^u[16]^u[14]^u[13]^u[11]^u[9]^u[8]^u[7]^u[6]^u[5]^u[3]^u[1]^u[0];
	y[174] = x[110]^x[237]^x[240]^x[242]^x[245]^x[247]^x[248]^x[249]^x[252]^x[254]^x[255]^x[257]^x[258]^x[259]^x[260]^x[266]^x[268]^x[272]^x[275]^x[281]^x[282]^x[284]^x[286]^x[287]^x[289]^x[291]^x[292]^x[293]^x[294]^x[295]^x[297]^x[299]^u[62]^u[59]^u[57]^u[54]^u[52]^u[51]^u[50]^u[47]^u[45]^u[44]^u[42]^u[41]^u[40]^u[39]^u[33]^u[31]^u[27]^u[24]^u[18]^u[17]^u[15]^u[13]^u[12]^u[10]^u[8]^u[7]^u[6]^u[5]^u[4]^u[2]^u[0];
	y[175] = x[111]^x[236]^x[239]^x[243]^x[245]^x[246]^x[248]^x[249]^x[250]^x[253]^x[256]^x[258]^x[259]^x[261]^x[264]^x[267]^x[271]^x[273]^x[279]^x[280]^x[282]^x[283]^x[288]^x[289]^x[290]^x[296]^u[63]^u[60]^u[56]^u[54]^u[53]^u[51]^u[50]^u[49]^u[46]^u[43]^u[41]^u[40]^u[38]^u[35]^u[32]^u[28]^u[26]^u[20]^u[19]^u[17]^u[16]^u[11]^u[10]^u[9]^u[3];
	y[176] = x[112]^x[237]^x[240]^x[244]^x[246]^x[247]^x[249]^x[250]^x[251]^x[254]^x[257]^x[259]^x[260]^x[262]^x[265]^x[268]^x[272]^x[274]^x[280]^x[281]^x[283]^x[284]^x[289]^x[290]^x[291]^x[297]^u[62]^u[59]^u[55]^u[53]^u[52]^u[50]^u[49]^u[48]^u[45]^u[42]^u[40]^u[39]^u[37]^u[34]^u[31]^u[27]^u[25]^u[19]^u[18]^u[16]^u[15]^u[10]^u[9]^u[8]^u[2];
	y[177] = x[113]^x[236]^x[239]^x[247]^x[248]^x[250]^x[251]^x[252]^x[258]^x[261]^x[263]^x[264]^x[266]^x[271]^x[273]^x[275]^x[276]^x[279]^x[280]^x[281]^x[282]^x[284]^x[287]^x[289]^x[290]^x[291]^x[293]^x[294]^x[295]^u[63]^u[60]^u[52]^u[51]^u[49]^u[48]^u[47]^u[41]^u[38]^u[36]^u[35]^u[33]^u[28]^u[26]^u[24]^u[23]^u[20]^u[19]^u[18]^u[17]^u[15]^u[12]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4];
	y[178] = x[114]^x[237]^x[240]^x[248]^x[249]^x[251]^x[252]^x[253]^x[259]^x[262]^x[264]^x[265]^x[267]^x[272]^x[274]^x[276]^x[277]^x[280]^x[281]^x[282]^x[283]^x[285]^x[288]^x[290]^x[291]^x[292]^x[294]^x[295]^x[296]^u[62]^u[59]^u[51]^u[50]^u[48]^u[47]^u[46]^u[40]^u[37]^u[35]^u[34]^u[32]^u[27]^u[25]^u[23]^u[22]^u[19]^u[18]^u[17]^u[16]^u[14]^u[11]^u[9]^u[8]^u[7]^u[5]^u[4]^u[3];
	y[179] = x[115]^x[238]^x[241]^x[249]^x[250]^x[252]^x[253]^x[254]^x[260]^x[263]^x[265]^x[266]^x[268]^x[273]^x[275]^x[277]^x[278]^x[281]^x[282]^x[283]^x[284]^x[286]^x[289]^x[291]^x[292]^x[293]^x[295]^x[296]^x[297]^u[61]^u[58]^u[50]^u[49]^u[47]^u[46]^u[45]^u[39]^u[36]^u[34]^u[33]^u[31]^u[26]^u[24]^u[22]^u[21]^u[18]^u[17]^u[16]^u[15]^u[13]^u[10]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2];
	y[180] = x[116]^x[239]^x[242]^x[250]^x[251]^x[253]^x[254]^x[255]^x[261]^x[264]^x[266]^x[267]^x[269]^x[274]^x[276]^x[278]^x[279]^x[282]^x[283]^x[284]^x[285]^x[287]^x[290]^x[292]^x[293]^x[294]^x[296]^x[297]^x[298]^u[60]^u[57]^u[49]^u[48]^u[46]^u[45]^u[44]^u[38]^u[35]^u[33]^u[32]^u[30]^u[25]^u[23]^u[21]^u[20]^u[17]^u[16]^u[15]^u[14]^u[12]^u[9]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[181] = x[117]^x[236]^x[238]^x[239]^x[240]^x[241]^x[243]^x[245]^x[251]^x[252]^x[254]^x[256]^x[260]^x[262]^x[264]^x[265]^x[267]^x[268]^x[269]^x[270]^x[271]^x[275]^x[276]^x[277]^x[283]^x[284]^x[286]^x[287]^x[288]^x[289]^x[291]^x[292]^x[297]^x[299]^u[63]^u[61]^u[60]^u[59]^u[58]^u[56]^u[54]^u[48]^u[47]^u[45]^u[43]^u[39]^u[37]^u[35]^u[34]^u[32]^u[31]^u[30]^u[29]^u[28]^u[24]^u[23]^u[22]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[8]^u[7]^u[2]^u[0];
	y[182] = x[118]^x[236]^x[237]^x[238]^x[240]^x[242]^x[244]^x[245]^x[246]^x[252]^x[253]^x[257]^x[260]^x[261]^x[263]^x[264]^x[265]^x[266]^x[268]^x[270]^x[272]^x[277]^x[278]^x[279]^x[280]^x[284]^x[288]^x[290]^x[294]^x[295]^u[63]^u[62]^u[61]^u[59]^u[57]^u[55]^u[54]^u[53]^u[47]^u[46]^u[42]^u[39]^u[38]^u[36]^u[35]^u[34]^u[33]^u[31]^u[29]^u[27]^u[22]^u[21]^u[20]^u[19]^u[15]^u[11]^u[9]^u[5]^u[4];
	y[183] = x[119]^x[237]^x[238]^x[239]^x[241]^x[243]^x[245]^x[246]^x[247]^x[253]^x[254]^x[258]^x[261]^x[262]^x[264]^x[265]^x[266]^x[267]^x[269]^x[271]^x[273]^x[278]^x[279]^x[280]^x[281]^x[285]^x[289]^x[291]^x[295]^x[296]^u[62]^u[61]^u[60]^u[58]^u[56]^u[54]^u[53]^u[52]^u[46]^u[45]^u[41]^u[38]^u[37]^u[35]^u[34]^u[33]^u[32]^u[30]^u[28]^u[26]^u[21]^u[20]^u[19]^u[18]^u[14]^u[10]^u[8]^u[4]^u[3];
	y[184] = x[120]^x[238]^x[239]^x[240]^x[242]^x[244]^x[246]^x[247]^x[248]^x[254]^x[255]^x[259]^x[262]^x[263]^x[265]^x[266]^x[267]^x[268]^x[270]^x[272]^x[274]^x[279]^x[280]^x[281]^x[282]^x[286]^x[290]^x[292]^x[296]^x[297]^u[61]^u[60]^u[59]^u[57]^u[55]^u[53]^u[52]^u[51]^u[45]^u[44]^u[40]^u[37]^u[36]^u[34]^u[33]^u[32]^u[31]^u[29]^u[27]^u[25]^u[20]^u[19]^u[18]^u[17]^u[13]^u[9]^u[7]^u[3]^u[2];
	y[185] = x[121]^x[239]^x[240]^x[241]^x[243]^x[245]^x[247]^x[248]^x[249]^x[255]^x[256]^x[260]^x[263]^x[264]^x[266]^x[267]^x[268]^x[269]^x[271]^x[273]^x[275]^x[280]^x[281]^x[282]^x[283]^x[287]^x[291]^x[293]^x[297]^x[298]^u[60]^u[59]^u[58]^u[56]^u[54]^u[52]^u[51]^u[50]^u[44]^u[43]^u[39]^u[36]^u[35]^u[33]^u[32]^u[31]^u[30]^u[28]^u[26]^u[24]^u[19]^u[18]^u[17]^u[16]^u[12]^u[8]^u[6]^u[2]^u[1];
	y[186] = x[122]^x[240]^x[241]^x[242]^x[244]^x[246]^x[248]^x[249]^x[250]^x[256]^x[257]^x[261]^x[264]^x[265]^x[267]^x[268]^x[269]^x[270]^x[272]^x[274]^x[276]^x[281]^x[282]^x[283]^x[284]^x[288]^x[292]^x[294]^x[298]^x[299]^u[59]^u[58]^u[57]^u[55]^u[53]^u[51]^u[50]^u[49]^u[43]^u[42]^u[38]^u[35]^u[34]^u[32]^u[31]^u[30]^u[29]^u[27]^u[25]^u[23]^u[18]^u[17]^u[16]^u[15]^u[11]^u[7]^u[5]^u[1]^u[0];
	y[187] = x[123]^x[236]^x[238]^x[239]^x[242]^x[243]^x[247]^x[249]^x[250]^x[251]^x[255]^x[257]^x[258]^x[260]^x[262]^x[264]^x[265]^x[266]^x[268]^x[270]^x[273]^x[275]^x[276]^x[277]^x[279]^x[280]^x[282]^x[283]^x[284]^x[287]^x[292]^x[294]^x[298]^x[299]^u[63]^u[61]^u[60]^u[57]^u[56]^u[52]^u[50]^u[49]^u[48]^u[44]^u[42]^u[41]^u[39]^u[37]^u[35]^u[34]^u[33]^u[31]^u[29]^u[26]^u[24]^u[23]^u[22]^u[20]^u[19]^u[17]^u[16]^u[15]^u[12]^u[7]^u[5]^u[1]^u[0];
	y[188] = x[124]^x[237]^x[239]^x[240]^x[243]^x[244]^x[248]^x[250]^x[251]^x[252]^x[256]^x[258]^x[259]^x[261]^x[263]^x[265]^x[266]^x[267]^x[269]^x[271]^x[274]^x[276]^x[277]^x[278]^x[280]^x[281]^x[283]^x[284]^x[285]^x[288]^x[293]^x[295]^x[299]^u[62]^u[60]^u[59]^u[56]^u[55]^u[51]^u[49]^u[48]^u[47]^u[43]^u[41]^u[40]^u[38]^u[36]^u[34]^u[33]^u[32]^u[30]^u[28]^u[25]^u[23]^u[22]^u[21]^u[19]^u[18]^u[16]^u[15]^u[14]^u[11]^u[6]^u[4]^u[0];
	y[189] = x[125]^x[238]^x[240]^x[241]^x[244]^x[245]^x[249]^x[251]^x[252]^x[253]^x[257]^x[259]^x[260]^x[262]^x[264]^x[266]^x[267]^x[268]^x[270]^x[272]^x[275]^x[277]^x[278]^x[279]^x[281]^x[282]^x[284]^x[285]^x[286]^x[289]^x[294]^x[296]^u[61]^u[59]^u[58]^u[55]^u[54]^u[50]^u[48]^u[47]^u[46]^u[42]^u[40]^u[39]^u[37]^u[35]^u[33]^u[32]^u[31]^u[29]^u[27]^u[24]^u[22]^u[21]^u[20]^u[18]^u[17]^u[15]^u[14]^u[13]^u[10]^u[5]^u[3];
	y[190] = x[126]^x[239]^x[241]^x[242]^x[245]^x[246]^x[250]^x[252]^x[253]^x[254]^x[258]^x[260]^x[261]^x[263]^x[265]^x[267]^x[268]^x[269]^x[271]^x[273]^x[276]^x[278]^x[279]^x[280]^x[282]^x[283]^x[285]^x[286]^x[287]^x[290]^x[295]^x[297]^u[60]^u[58]^u[57]^u[54]^u[53]^u[49]^u[47]^u[46]^u[45]^u[41]^u[39]^u[38]^u[36]^u[34]^u[32]^u[31]^u[30]^u[28]^u[26]^u[23]^u[21]^u[20]^u[19]^u[17]^u[16]^u[14]^u[13]^u[12]^u[9]^u[4]^u[2];
	y[191] = x[127]^x[240]^x[242]^x[243]^x[246]^x[247]^x[251]^x[253]^x[254]^x[255]^x[259]^x[261]^x[262]^x[264]^x[266]^x[268]^x[269]^x[270]^x[272]^x[274]^x[277]^x[279]^x[280]^x[281]^x[283]^x[284]^x[286]^x[287]^x[288]^x[291]^x[296]^x[298]^u[59]^u[57]^u[56]^u[53]^u[52]^u[48]^u[46]^u[45]^u[44]^u[40]^u[38]^u[37]^u[35]^u[33]^u[31]^u[30]^u[29]^u[27]^u[25]^u[22]^u[20]^u[19]^u[18]^u[16]^u[15]^u[13]^u[12]^u[11]^u[8]^u[3]^u[1];
	y[192] = x[128]^x[236]^x[238]^x[239]^x[243]^x[244]^x[245]^x[247]^x[248]^x[252]^x[254]^x[256]^x[262]^x[263]^x[264]^x[265]^x[267]^x[270]^x[273]^x[275]^x[276]^x[278]^x[279]^x[281]^x[282]^x[284]^x[288]^x[293]^x[294]^x[295]^x[297]^x[298]^x[299]^u[63]^u[61]^u[60]^u[56]^u[55]^u[54]^u[52]^u[51]^u[47]^u[45]^u[43]^u[37]^u[36]^u[35]^u[34]^u[32]^u[29]^u[26]^u[24]^u[23]^u[21]^u[20]^u[18]^u[17]^u[15]^u[11]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[193] = x[129]^x[236]^x[237]^x[238]^x[240]^x[241]^x[244]^x[246]^x[248]^x[249]^x[253]^x[257]^x[260]^x[263]^x[265]^x[266]^x[268]^x[269]^x[274]^x[277]^x[282]^x[283]^x[287]^x[292]^x[293]^x[296]^x[299]^u[63]^u[62]^u[61]^u[59]^u[58]^u[55]^u[53]^u[51]^u[50]^u[46]^u[42]^u[39]^u[36]^u[34]^u[33]^u[31]^u[30]^u[25]^u[22]^u[17]^u[16]^u[12]^u[7]^u[6]^u[3]^u[0];
	y[194] = x[130]^x[236]^x[237]^x[242]^x[247]^x[249]^x[250]^x[254]^x[255]^x[258]^x[260]^x[261]^x[266]^x[267]^x[270]^x[271]^x[275]^x[276]^x[278]^x[279]^x[280]^x[283]^x[284]^x[285]^x[287]^x[288]^x[289]^x[292]^x[295]^x[297]^x[298]^u[63]^u[62]^u[57]^u[52]^u[50]^u[49]^u[45]^u[44]^u[41]^u[39]^u[38]^u[33]^u[32]^u[29]^u[28]^u[24]^u[23]^u[21]^u[20]^u[19]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[7]^u[4]^u[2]^u[1];
	y[195] = x[131]^x[237]^x[238]^x[243]^x[248]^x[250]^x[251]^x[255]^x[256]^x[259]^x[261]^x[262]^x[267]^x[268]^x[271]^x[272]^x[276]^x[277]^x[279]^x[280]^x[281]^x[284]^x[285]^x[286]^x[288]^x[289]^x[290]^x[293]^x[296]^x[298]^x[299]^u[62]^u[61]^u[56]^u[51]^u[49]^u[48]^u[44]^u[43]^u[40]^u[38]^u[37]^u[32]^u[31]^u[28]^u[27]^u[23]^u[22]^u[20]^u[19]^u[18]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[6]^u[3]^u[1]^u[0];
	y[196] = x[132]^x[238]^x[239]^x[244]^x[249]^x[251]^x[252]^x[256]^x[257]^x[260]^x[262]^x[263]^x[268]^x[269]^x[272]^x[273]^x[277]^x[278]^x[280]^x[281]^x[282]^x[285]^x[286]^x[287]^x[289]^x[290]^x[291]^x[294]^x[297]^x[299]^u[61]^u[60]^u[55]^u[50]^u[48]^u[47]^u[43]^u[42]^u[39]^u[37]^u[36]^u[31]^u[30]^u[27]^u[26]^u[22]^u[21]^u[19]^u[18]^u[17]^u[14]^u[13]^u[12]^u[10]^u[9]^u[8]^u[5]^u[2]^u[0];
	y[197] = x[133]^x[236]^x[238]^x[240]^x[241]^x[250]^x[252]^x[253]^x[255]^x[257]^x[258]^x[260]^x[261]^x[263]^x[270]^x[271]^x[273]^x[274]^x[276]^x[278]^x[280]^x[281]^x[282]^x[283]^x[285]^x[286]^x[288]^x[289]^x[290]^x[291]^x[293]^x[294]^u[63]^u[61]^u[59]^u[58]^u[49]^u[47]^u[46]^u[44]^u[42]^u[41]^u[39]^u[38]^u[36]^u[29]^u[28]^u[26]^u[25]^u[23]^u[21]^u[19]^u[18]^u[17]^u[16]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[6]^u[5];
	y[198] = x[134]^x[237]^x[239]^x[241]^x[242]^x[251]^x[253]^x[254]^x[256]^x[258]^x[259]^x[261]^x[262]^x[264]^x[271]^x[272]^x[274]^x[275]^x[277]^x[279]^x[281]^x[282]^x[283]^x[284]^x[286]^x[287]^x[289]^x[290]^x[291]^x[292]^x[294]^x[295]^u[62]^u[60]^u[58]^u[57]^u[48]^u[46]^u[45]^u[43]^u[41]^u[40]^u[38]^u[37]^u[35]^u[28]^u[27]^u[25]^u[24]^u[22]^u[20]^u[18]^u[17]^u[16]^u[15]^u[13]^u[12]^u[10]^u[9]^u[8]^u[7]^u[5]^u[4];
	y[199] = x[135]^x[238]^x[240]^x[242]^x[243]^x[252]^x[254]^x[255]^x[257]^x[259]^x[260]^x[262]^x[263]^x[265]^x[272]^x[273]^x[275]^x[276]^x[278]^x[280]^x[282]^x[283]^x[284]^x[285]^x[287]^x[288]^x[290]^x[291]^x[292]^x[293]^x[295]^x[296]^u[61]^u[59]^u[57]^u[56]^u[47]^u[45]^u[44]^u[42]^u[40]^u[39]^u[37]^u[36]^u[34]^u[27]^u[26]^u[24]^u[23]^u[21]^u[19]^u[17]^u[16]^u[15]^u[14]^u[12]^u[11]^u[9]^u[8]^u[7]^u[6]^u[4]^u[3];
	y[200] = x[136]^x[239]^x[241]^x[243]^x[244]^x[253]^x[255]^x[256]^x[258]^x[260]^x[261]^x[263]^x[264]^x[266]^x[273]^x[274]^x[276]^x[277]^x[279]^x[281]^x[283]^x[284]^x[285]^x[286]^x[288]^x[289]^x[291]^x[292]^x[293]^x[294]^x[296]^x[297]^u[60]^u[58]^u[56]^u[55]^u[46]^u[44]^u[43]^u[41]^u[39]^u[38]^u[36]^u[35]^u[33]^u[26]^u[25]^u[23]^u[22]^u[20]^u[18]^u[16]^u[15]^u[14]^u[13]^u[11]^u[10]^u[8]^u[7]^u[6]^u[5]^u[3]^u[2];
	y[201] = x[137]^x[240]^x[242]^x[244]^x[245]^x[254]^x[256]^x[257]^x[259]^x[261]^x[262]^x[264]^x[265]^x[267]^x[274]^x[275]^x[277]^x[278]^x[280]^x[282]^x[284]^x[285]^x[286]^x[287]^x[289]^x[290]^x[292]^x[293]^x[294]^x[295]^x[297]^x[298]^u[59]^u[57]^u[55]^u[54]^u[45]^u[43]^u[42]^u[40]^u[38]^u[37]^u[35]^u[34]^u[32]^u[25]^u[24]^u[22]^u[21]^u[19]^u[17]^u[15]^u[14]^u[13]^u[12]^u[10]^u[9]^u[7]^u[6]^u[5]^u[4]^u[2]^u[1];
	y[202] = x[138]^x[236]^x[238]^x[239]^x[243]^x[246]^x[257]^x[258]^x[262]^x[263]^x[264]^x[265]^x[266]^x[268]^x[269]^x[271]^x[275]^x[278]^x[280]^x[281]^x[283]^x[286]^x[288]^x[289]^x[290]^x[291]^x[292]^x[296]^x[299]^u[63]^u[61]^u[60]^u[56]^u[53]^u[42]^u[41]^u[37]^u[36]^u[35]^u[34]^u[33]^u[31]^u[30]^u[28]^u[24]^u[21]^u[19]^u[18]^u[16]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[3]^u[0];
	y[203] = x[139]^x[236]^x[237]^x[238]^x[240]^x[241]^x[244]^x[245]^x[247]^x[255]^x[258]^x[259]^x[260]^x[263]^x[265]^x[266]^x[267]^x[270]^x[271]^x[272]^x[280]^x[281]^x[282]^x[284]^x[285]^x[290]^x[291]^x[294]^x[295]^x[297]^x[298]^u[63]^u[62]^u[61]^u[59]^u[58]^u[55]^u[54]^u[52]^u[44]^u[41]^u[40]^u[39]^u[36]^u[34]^u[33]^u[32]^u[29]^u[28]^u[27]^u[19]^u[18]^u[17]^u[15]^u[14]^u[9]^u[8]^u[5]^u[4]^u[2]^u[1];
	y[204] = x[140]^x[236]^x[237]^x[242]^x[246]^x[248]^x[255]^x[256]^x[259]^x[261]^x[266]^x[267]^x[268]^x[269]^x[272]^x[273]^x[276]^x[279]^x[280]^x[281]^x[282]^x[283]^x[286]^x[287]^x[289]^x[291]^x[293]^x[294]^x[296]^x[299]^u[63]^u[62]^u[57]^u[53]^u[51]^u[44]^u[43]^u[40]^u[38]^u[33]^u[32]^u[31]^u[30]^u[27]^u[26]^u[23]^u[20]^u[19]^u[18]^u[17]^u[16]^u[13]^u[12]^u[10]^u[8]^u[6]^u[5]^u[3]^u[0];
	y[205] = x[141]^x[237]^x[238]^x[243]^x[247]^x[249]^x[256]^x[257]^x[260]^x[262]^x[267]^x[268]^x[269]^x[270]^x[273]^x[274]^x[277]^x[280]^x[281]^x[282]^x[283]^x[284]^x[287]^x[288]^x[290]^x[292]^x[294]^x[295]^x[297]^u[62]^u[61]^u[56]^u[52]^u[50]^u[43]^u[42]^u[39]^u[37]^u[32]^u[31]^u[30]^u[29]^u[26]^u[25]^u[22]^u[19]^u[18]^u[17]^u[16]^u[15]^u[12]^u[11]^u[9]^u[7]^u[5]^u[4]^u[2];
	y[206] = x[142]^x[238]^x[239]^x[244]^x[248]^x[250]^x[257]^x[258]^x[261]^x[263]^x[268]^x[269]^x[270]^x[271]^x[274]^x[275]^x[278]^x[281]^x[282]^x[283]^x[284]^x[285]^x[288]^x[289]^x[291]^x[293]^x[295]^x[296]^x[298]^u[61]^u[60]^u[55]^u[51]^u[49]^u[42]^u[41]^u[38]^u[36]^u[31]^u[30]^u[29]^u[28]^u[25]^u[24]^u[21]^u[18]^u[17]^u[16]^u[15]^u[14]^u[11]^u[10]^u[8]^u[6]^u[4]^u[3]^u[1];
	y[207] = x[143]^x[236]^x[238]^x[240]^x[241]^x[249]^x[251]^x[255]^x[258]^x[259]^x[260]^x[262]^x[270]^x[272]^x[275]^x[280]^x[282]^x[283]^x[284]^x[286]^x[287]^x[290]^x[293]^x[295]^x[296]^x[297]^x[298]^x[299]^u[63]^u[61]^u[59]^u[58]^u[50]^u[48]^u[44]^u[41]^u[40]^u[39]^u[37]^u[29]^u[27]^u[24]^u[19]^u[17]^u[16]^u[15]^u[13]^u[12]^u[9]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[208] = x[144]^x[236]^x[237]^x[238]^x[242]^x[245]^x[250]^x[252]^x[255]^x[256]^x[259]^x[261]^x[263]^x[264]^x[269]^x[273]^x[279]^x[280]^x[281]^x[283]^x[284]^x[288]^x[289]^x[291]^x[292]^x[293]^x[295]^x[296]^x[297]^x[299]^u[63]^u[62]^u[61]^u[57]^u[54]^u[49]^u[47]^u[44]^u[43]^u[40]^u[38]^u[36]^u[35]^u[30]^u[26]^u[20]^u[19]^u[18]^u[16]^u[15]^u[11]^u[10]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[0];
	y[209] = x[145]^x[237]^x[238]^x[239]^x[243]^x[246]^x[251]^x[253]^x[256]^x[257]^x[260]^x[262]^x[264]^x[265]^x[270]^x[274]^x[280]^x[281]^x[282]^x[284]^x[285]^x[289]^x[290]^x[292]^x[293]^x[294]^x[296]^x[297]^x[298]^u[62]^u[61]^u[60]^u[56]^u[53]^u[48]^u[46]^u[43]^u[42]^u[39]^u[37]^u[35]^u[34]^u[29]^u[25]^u[19]^u[18]^u[17]^u[15]^u[14]^u[10]^u[9]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[210] = x[146]^x[238]^x[239]^x[240]^x[244]^x[247]^x[252]^x[254]^x[257]^x[258]^x[261]^x[263]^x[265]^x[266]^x[271]^x[275]^x[281]^x[282]^x[283]^x[285]^x[286]^x[290]^x[291]^x[293]^x[294]^x[295]^x[297]^x[298]^x[299]^u[61]^u[60]^u[59]^u[55]^u[52]^u[47]^u[45]^u[42]^u[41]^u[38]^u[36]^u[34]^u[33]^u[28]^u[24]^u[18]^u[17]^u[16]^u[14]^u[13]^u[9]^u[8]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[211] = x[147]^x[239]^x[240]^x[241]^x[245]^x[248]^x[253]^x[255]^x[258]^x[259]^x[262]^x[264]^x[266]^x[267]^x[272]^x[276]^x[282]^x[283]^x[284]^x[286]^x[287]^x[291]^x[292]^x[294]^x[295]^x[296]^x[298]^x[299]^u[60]^u[59]^u[58]^u[54]^u[51]^u[46]^u[44]^u[41]^u[40]^u[37]^u[35]^u[33]^u[32]^u[27]^u[23]^u[17]^u[16]^u[15]^u[13]^u[12]^u[8]^u[7]^u[5]^u[4]^u[3]^u[1]^u[0];
	y[212] = x[148]^x[240]^x[241]^x[242]^x[246]^x[249]^x[254]^x[256]^x[259]^x[260]^x[263]^x[265]^x[267]^x[268]^x[273]^x[277]^x[283]^x[284]^x[285]^x[287]^x[288]^x[292]^x[293]^x[295]^x[296]^x[297]^x[299]^u[59]^u[58]^u[57]^u[53]^u[50]^u[45]^u[43]^u[40]^u[39]^u[36]^u[34]^u[32]^u[31]^u[26]^u[22]^u[16]^u[15]^u[14]^u[12]^u[11]^u[7]^u[6]^u[4]^u[3]^u[2]^u[0];
	y[213] = x[149]^x[241]^x[242]^x[243]^x[247]^x[250]^x[255]^x[257]^x[260]^x[261]^x[264]^x[266]^x[268]^x[269]^x[274]^x[278]^x[284]^x[285]^x[286]^x[288]^x[289]^x[293]^x[294]^x[296]^x[297]^x[298]^u[58]^u[57]^u[56]^u[52]^u[49]^u[44]^u[42]^u[39]^u[38]^u[35]^u[33]^u[31]^u[30]^u[25]^u[21]^u[15]^u[14]^u[13]^u[11]^u[10]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[214] = x[150]^x[236]^x[238]^x[239]^x[241]^x[242]^x[243]^x[244]^x[245]^x[248]^x[251]^x[255]^x[256]^x[258]^x[260]^x[261]^x[262]^x[264]^x[265]^x[267]^x[270]^x[271]^x[275]^x[276]^x[280]^x[286]^x[290]^x[292]^x[293]^x[297]^x[299]^u[63]^u[61]^u[60]^u[58]^u[57]^u[56]^u[55]^u[54]^u[51]^u[48]^u[44]^u[43]^u[41]^u[39]^u[38]^u[37]^u[35]^u[34]^u[32]^u[29]^u[28]^u[24]^u[23]^u[19]^u[13]^u[9]^u[7]^u[6]^u[2]^u[0];
	y[215] = x[151]^x[237]^x[239]^x[240]^x[242]^x[243]^x[244]^x[245]^x[246]^x[249]^x[252]^x[256]^x[257]^x[259]^x[261]^x[262]^x[263]^x[265]^x[266]^x[268]^x[271]^x[272]^x[276]^x[277]^x[281]^x[287]^x[291]^x[293]^x[294]^x[298]^u[62]^u[60]^u[59]^u[57]^u[56]^u[55]^u[54]^u[53]^u[50]^u[47]^u[43]^u[42]^u[40]^u[38]^u[37]^u[36]^u[34]^u[33]^u[31]^u[28]^u[27]^u[23]^u[22]^u[18]^u[12]^u[8]^u[6]^u[5]^u[1];
	y[216] = x[152]^x[238]^x[240]^x[241]^x[243]^x[244]^x[245]^x[246]^x[247]^x[250]^x[253]^x[257]^x[258]^x[260]^x[262]^x[263]^x[264]^x[266]^x[267]^x[269]^x[272]^x[273]^x[277]^x[278]^x[282]^x[288]^x[292]^x[294]^x[295]^x[299]^u[61]^u[59]^u[58]^u[56]^u[55]^u[54]^u[53]^u[52]^u[49]^u[46]^u[42]^u[41]^u[39]^u[37]^u[36]^u[35]^u[33]^u[32]^u[30]^u[27]^u[26]^u[22]^u[21]^u[17]^u[11]^u[7]^u[5]^u[4]^u[0];
	y[217] = x[153]^x[236]^x[238]^x[242]^x[244]^x[246]^x[247]^x[248]^x[251]^x[254]^x[255]^x[258]^x[259]^x[260]^x[261]^x[263]^x[265]^x[267]^x[268]^x[269]^x[270]^x[271]^x[273]^x[274]^x[276]^x[278]^x[280]^x[283]^x[285]^x[287]^x[292]^x[294]^x[296]^x[298]^u[63]^u[61]^u[57]^u[55]^u[53]^u[52]^u[51]^u[48]^u[45]^u[44]^u[41]^u[40]^u[39]^u[38]^u[36]^u[34]^u[32]^u[31]^u[30]^u[29]^u[28]^u[26]^u[25]^u[23]^u[21]^u[19]^u[16]^u[14]^u[12]^u[7]^u[5]^u[3]^u[1];
	y[218] = x[154]^x[237]^x[239]^x[243]^x[245]^x[247]^x[248]^x[249]^x[252]^x[255]^x[256]^x[259]^x[260]^x[261]^x[262]^x[264]^x[266]^x[268]^x[269]^x[270]^x[271]^x[272]^x[274]^x[275]^x[277]^x[279]^x[281]^x[284]^x[286]^x[288]^x[293]^x[295]^x[297]^x[299]^u[62]^u[60]^u[56]^u[54]^u[52]^u[51]^u[50]^u[47]^u[44]^u[43]^u[40]^u[39]^u[38]^u[37]^u[35]^u[33]^u[31]^u[30]^u[29]^u[28]^u[27]^u[25]^u[24]^u[22]^u[20]^u[18]^u[15]^u[13]^u[11]^u[6]^u[4]^u[2]^u[0];
	y[219] = x[155]^x[236]^x[239]^x[240]^x[241]^x[244]^x[245]^x[246]^x[248]^x[249]^x[250]^x[253]^x[255]^x[256]^x[257]^x[261]^x[262]^x[263]^x[264]^x[265]^x[267]^x[270]^x[272]^x[273]^x[275]^x[278]^x[279]^x[282]^x[292]^x[293]^x[295]^x[296]^u[63]^u[60]^u[59]^u[58]^u[55]^u[54]^u[53]^u[51]^u[50]^u[49]^u[46]^u[44]^u[43]^u[42]^u[38]^u[37]^u[36]^u[35]^u[34]^u[32]^u[29]^u[27]^u[26]^u[24]^u[21]^u[20]^u[17]^u[7]^u[6]^u[4]^u[3];
	y[220] = x[156]^x[237]^x[240]^x[241]^x[242]^x[245]^x[246]^x[247]^x[249]^x[250]^x[251]^x[254]^x[256]^x[257]^x[258]^x[262]^x[263]^x[264]^x[265]^x[266]^x[268]^x[271]^x[273]^x[274]^x[276]^x[279]^x[280]^x[283]^x[293]^x[294]^x[296]^x[297]^u[62]^u[59]^u[58]^u[57]^u[54]^u[53]^u[52]^u[50]^u[49]^u[48]^u[45]^u[43]^u[42]^u[41]^u[37]^u[36]^u[35]^u[34]^u[33]^u[31]^u[28]^u[26]^u[25]^u[23]^u[20]^u[19]^u[16]^u[6]^u[5]^u[3]^u[2];
	y[221] = x[157]^x[238]^x[241]^x[242]^x[243]^x[246]^x[247]^x[248]^x[250]^x[251]^x[252]^x[255]^x[257]^x[258]^x[259]^x[263]^x[264]^x[265]^x[266]^x[267]^x[269]^x[272]^x[274]^x[275]^x[277]^x[280]^x[281]^x[284]^x[294]^x[295]^x[297]^x[298]^u[61]^u[58]^u[57]^u[56]^u[53]^u[52]^u[51]^u[49]^u[48]^u[47]^u[44]^u[42]^u[41]^u[40]^u[36]^u[35]^u[34]^u[33]^u[32]^u[30]^u[27]^u[25]^u[24]^u[22]^u[19]^u[18]^u[15]^u[5]^u[4]^u[2]^u[1];
	y[222] = x[158]^x[236]^x[238]^x[241]^x[242]^x[243]^x[244]^x[245]^x[247]^x[248]^x[249]^x[251]^x[252]^x[253]^x[255]^x[256]^x[258]^x[259]^x[265]^x[266]^x[267]^x[268]^x[269]^x[270]^x[271]^x[273]^x[275]^x[278]^x[279]^x[280]^x[281]^x[282]^x[287]^x[289]^x[292]^x[293]^x[294]^x[296]^x[299]^u[63]^u[61]^u[58]^u[57]^u[56]^u[55]^u[54]^u[52]^u[51]^u[50]^u[48]^u[47]^u[46]^u[44]^u[43]^u[41]^u[40]^u[34]^u[33]^u[32]^u[31]^u[30]^u[29]^u[28]^u[26]^u[24]^u[21]^u[20]^u[19]^u[18]^u[17]^u[12]^u[10]^u[7]^u[6]^u[5]^u[3]^u[0];
	y[223] = x[159]^x[236]^x[237]^x[238]^x[241]^x[242]^x[243]^x[244]^x[246]^x[248]^x[249]^x[250]^x[252]^x[253]^x[254]^x[255]^x[256]^x[257]^x[259]^x[264]^x[266]^x[267]^x[268]^x[270]^x[272]^x[274]^x[281]^x[282]^x[283]^x[285]^x[287]^x[288]^x[289]^x[290]^x[292]^x[297]^x[298]^u[63]^u[62]^u[61]^u[58]^u[57]^u[56]^u[55]^u[53]^u[51]^u[50]^u[49]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[40]^u[35]^u[33]^u[32]^u[31]^u[29]^u[27]^u[25]^u[18]^u[17]^u[16]^u[14]^u[12]^u[11]^u[10]^u[9]^u[7]^u[2]^u[1];
	y[224] = x[160]^x[236]^x[237]^x[241]^x[242]^x[243]^x[244]^x[247]^x[249]^x[250]^x[251]^x[253]^x[254]^x[256]^x[257]^x[258]^x[264]^x[265]^x[267]^x[268]^x[273]^x[275]^x[276]^x[279]^x[280]^x[282]^x[283]^x[284]^x[285]^x[286]^x[287]^x[288]^x[290]^x[291]^x[292]^x[294]^x[295]^x[299]^u[63]^u[62]^u[58]^u[57]^u[56]^u[55]^u[52]^u[50]^u[49]^u[48]^u[46]^u[45]^u[43]^u[42]^u[41]^u[35]^u[34]^u[32]^u[31]^u[26]^u[24]^u[23]^u[20]^u[19]^u[17]^u[16]^u[15]^u[14]^u[13]^u[12]^u[11]^u[9]^u[8]^u[7]^u[5]^u[4]^u[0];
	y[225] = x[161]^x[236]^x[237]^x[239]^x[241]^x[242]^x[243]^x[244]^x[248]^x[250]^x[251]^x[252]^x[254]^x[257]^x[258]^x[259]^x[260]^x[264]^x[265]^x[266]^x[268]^x[271]^x[274]^x[277]^x[279]^x[281]^x[283]^x[284]^x[286]^x[288]^x[291]^x[294]^x[296]^x[298]^u[63]^u[62]^u[60]^u[58]^u[57]^u[56]^u[55]^u[51]^u[49]^u[48]^u[47]^u[45]^u[42]^u[41]^u[40]^u[39]^u[35]^u[34]^u[33]^u[31]^u[28]^u[25]^u[22]^u[20]^u[18]^u[16]^u[15]^u[13]^u[11]^u[8]^u[5]^u[3]^u[1];
	y[226] = x[162]^x[236]^x[237]^x[239]^x[240]^x[241]^x[242]^x[243]^x[244]^x[249]^x[251]^x[252]^x[253]^x[258]^x[259]^x[261]^x[264]^x[265]^x[266]^x[267]^x[271]^x[272]^x[275]^x[276]^x[278]^x[279]^x[282]^x[284]^x[293]^x[294]^x[297]^x[298]^x[299]^u[63]^u[62]^u[60]^u[59]^u[58]^u[57]^u[56]^u[55]^u[50]^u[48]^u[47]^u[46]^u[41]^u[40]^u[38]^u[35]^u[34]^u[33]^u[32]^u[28]^u[27]^u[24]^u[23]^u[21]^u[20]^u[17]^u[15]^u[6]^u[5]^u[2]^u[1]^u[0];
	y[227] = x[163]^x[237]^x[238]^x[240]^x[241]^x[242]^x[243]^x[244]^x[245]^x[250]^x[252]^x[253]^x[254]^x[259]^x[260]^x[262]^x[265]^x[266]^x[267]^x[268]^x[272]^x[273]^x[276]^x[277]^x[279]^x[280]^x[283]^x[285]^x[294]^x[295]^x[298]^x[299]^u[62]^u[61]^u[59]^u[58]^u[57]^u[56]^u[55]^u[54]^u[49]^u[47]^u[46]^u[45]^u[40]^u[39]^u[37]^u[34]^u[33]^u[32]^u[31]^u[27]^u[26]^u[23]^u[22]^u[20]^u[19]^u[16]^u[14]^u[5]^u[4]^u[1]^u[0];
	y[228] = x[164]^x[236]^x[242]^x[243]^x[244]^x[246]^x[251]^x[253]^x[254]^x[261]^x[263]^x[264]^x[266]^x[267]^x[268]^x[271]^x[273]^x[274]^x[276]^x[277]^x[278]^x[279]^x[281]^x[284]^x[285]^x[286]^x[287]^x[289]^x[292]^x[293]^x[294]^x[296]^x[298]^x[299]^u[63]^u[57]^u[56]^u[55]^u[53]^u[48]^u[46]^u[45]^u[38]^u[36]^u[35]^u[33]^u[32]^u[31]^u[28]^u[26]^u[25]^u[23]^u[22]^u[21]^u[20]^u[18]^u[15]^u[14]^u[13]^u[12]^u[10]^u[7]^u[6]^u[5]^u[3]^u[1]^u[0];
	y[229] = x[165]^x[236]^x[237]^x[238]^x[239]^x[241]^x[243]^x[244]^x[247]^x[252]^x[254]^x[260]^x[262]^x[265]^x[267]^x[268]^x[271]^x[272]^x[274]^x[275]^x[276]^x[277]^x[278]^x[282]^x[286]^x[288]^x[289]^x[290]^x[292]^x[297]^x[298]^x[299]^u[63]^u[62]^u[61]^u[60]^u[58]^u[56]^u[55]^u[52]^u[47]^u[45]^u[39]^u[37]^u[34]^u[32]^u[31]^u[28]^u[27]^u[25]^u[24]^u[23]^u[22]^u[21]^u[17]^u[13]^u[11]^u[10]^u[9]^u[7]^u[2]^u[1]^u[0];
	y[230] = x[166]^x[237]^x[238]^x[239]^x[240]^x[242]^x[244]^x[245]^x[248]^x[253]^x[255]^x[261]^x[263]^x[266]^x[268]^x[269]^x[272]^x[273]^x[275]^x[276]^x[277]^x[278]^x[279]^x[283]^x[287]^x[289]^x[290]^x[291]^x[293]^x[298]^x[299]^u[62]^u[61]^u[60]^u[59]^u[57]^u[55]^u[54]^u[51]^u[46]^u[44]^u[38]^u[36]^u[33]^u[31]^u[30]^u[27]^u[26]^u[24]^u[23]^u[22]^u[21]^u[20]^u[16]^u[12]^u[10]^u[9]^u[8]^u[6]^u[1]^u[0];
	y[231] = x[167]^x[238]^x[239]^x[240]^x[241]^x[243]^x[245]^x[246]^x[249]^x[254]^x[256]^x[262]^x[264]^x[267]^x[269]^x[270]^x[273]^x[274]^x[276]^x[277]^x[278]^x[279]^x[280]^x[284]^x[288]^x[290]^x[291]^x[292]^x[294]^x[299]^u[61]^u[60]^u[59]^u[58]^u[56]^u[54]^u[53]^u[50]^u[45]^u[43]^u[37]^u[35]^u[32]^u[30]^u[29]^u[26]^u[25]^u[23]^u[22]^u[21]^u[20]^u[19]^u[15]^u[11]^u[9]^u[8]^u[7]^u[5]^u[0];
	y[232] = x[168]^x[239]^x[240]^x[241]^x[242]^x[244]^x[246]^x[247]^x[250]^x[255]^x[257]^x[263]^x[265]^x[268]^x[270]^x[271]^x[274]^x[275]^x[277]^x[278]^x[279]^x[280]^x[281]^x[285]^x[289]^x[291]^x[292]^x[293]^x[295]^u[60]^u[59]^u[58]^u[57]^u[55]^u[53]^u[52]^u[49]^u[44]^u[42]^u[36]^u[34]^u[31]^u[29]^u[28]^u[25]^u[24]^u[22]^u[21]^u[20]^u[19]^u[18]^u[14]^u[10]^u[8]^u[7]^u[6]^u[4];
	y[233] = x[169]^x[236]^x[238]^x[239]^x[240]^x[242]^x[243]^x[247]^x[248]^x[251]^x[255]^x[256]^x[258]^x[260]^x[266]^x[272]^x[275]^x[278]^x[281]^x[282]^x[285]^x[286]^x[287]^x[289]^x[290]^x[295]^x[296]^x[298]^u[63]^u[61]^u[60]^u[59]^u[57]^u[56]^u[52]^u[51]^u[48]^u[44]^u[43]^u[41]^u[39]^u[33]^u[27]^u[24]^u[21]^u[18]^u[17]^u[14]^u[13]^u[12]^u[10]^u[9]^u[4]^u[3]^u[1];
	y[234] = x[170]^x[237]^x[239]^x[240]^x[241]^x[243]^x[244]^x[248]^x[249]^x[252]^x[256]^x[257]^x[259]^x[261]^x[267]^x[273]^x[276]^x[279]^x[282]^x[283]^x[286]^x[287]^x[288]^x[290]^x[291]^x[296]^x[297]^x[299]^u[62]^u[60]^u[59]^u[58]^u[56]^u[55]^u[51]^u[50]^u[47]^u[43]^u[42]^u[40]^u[38]^u[32]^u[26]^u[23]^u[20]^u[17]^u[16]^u[13]^u[12]^u[11]^u[9]^u[8]^u[3]^u[2]^u[0];
	y[235] = x[171]^x[236]^x[239]^x[240]^x[242]^x[244]^x[249]^x[250]^x[253]^x[255]^x[257]^x[258]^x[262]^x[264]^x[268]^x[269]^x[271]^x[274]^x[276]^x[277]^x[279]^x[283]^x[284]^x[285]^x[288]^x[291]^x[293]^x[294]^x[295]^x[297]^u[63]^u[60]^u[59]^u[57]^u[55]^u[50]^u[49]^u[46]^u[44]^u[42]^u[41]^u[37]^u[35]^u[31]^u[30]^u[28]^u[25]^u[23]^u[22]^u[20]^u[16]^u[15]^u[14]^u[11]^u[8]^u[6]^u[5]^u[4]^u[2];
	y[236] = x[172]^x[237]^x[240]^x[241]^x[243]^x[245]^x[250]^x[251]^x[254]^x[256]^x[258]^x[259]^x[263]^x[265]^x[269]^x[270]^x[272]^x[275]^x[277]^x[278]^x[280]^x[284]^x[285]^x[286]^x[289]^x[292]^x[294]^x[295]^x[296]^x[298]^u[62]^u[59]^u[58]^u[56]^u[54]^u[49]^u[48]^u[45]^u[43]^u[41]^u[40]^u[36]^u[34]^u[30]^u[29]^u[27]^u[24]^u[22]^u[21]^u[19]^u[15]^u[14]^u[13]^u[10]^u[7]^u[5]^u[4]^u[3]^u[1];
	y[237] = x[173]^x[236]^x[239]^x[242]^x[244]^x[245]^x[246]^x[251]^x[252]^x[257]^x[259]^x[266]^x[269]^x[270]^x[273]^x[278]^x[280]^x[281]^x[286]^x[289]^x[290]^x[292]^x[294]^x[296]^x[297]^x[298]^x[299]^u[63]^u[60]^u[57]^u[55]^u[54]^u[53]^u[48]^u[47]^u[42]^u[40]^u[33]^u[30]^u[29]^u[26]^u[21]^u[19]^u[18]^u[13]^u[10]^u[9]^u[7]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[238] = x[174]^x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[243]^x[246]^x[247]^x[252]^x[253]^x[255]^x[258]^x[264]^x[267]^x[269]^x[270]^x[274]^x[276]^x[280]^x[281]^x[282]^x[285]^x[289]^x[290]^x[291]^x[292]^x[294]^x[297]^x[299]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[56]^u[53]^u[52]^u[47]^u[46]^u[44]^u[41]^u[35]^u[32]^u[30]^u[29]^u[25]^u[23]^u[19]^u[18]^u[17]^u[14]^u[10]^u[9]^u[8]^u[7]^u[5]^u[2]^u[0];
	y[239] = x[175]^x[237]^x[238]^x[239]^x[240]^x[241]^x[242]^x[244]^x[247]^x[248]^x[253]^x[254]^x[256]^x[259]^x[265]^x[268]^x[270]^x[271]^x[275]^x[277]^x[281]^x[282]^x[283]^x[286]^x[290]^x[291]^x[292]^x[293]^x[295]^x[298]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[55]^u[52]^u[51]^u[46]^u[45]^u[43]^u[40]^u[34]^u[31]^u[29]^u[28]^u[24]^u[22]^u[18]^u[17]^u[16]^u[13]^u[9]^u[8]^u[7]^u[6]^u[4]^u[1];
	y[240] = x[176]^x[238]^x[239]^x[240]^x[241]^x[242]^x[243]^x[245]^x[248]^x[249]^x[254]^x[255]^x[257]^x[260]^x[266]^x[269]^x[271]^x[272]^x[276]^x[278]^x[282]^x[283]^x[284]^x[287]^x[291]^x[292]^x[293]^x[294]^x[296]^x[299]^u[61]^u[60]^u[59]^u[58]^u[57]^u[56]^u[54]^u[51]^u[50]^u[45]^u[44]^u[42]^u[39]^u[33]^u[30]^u[28]^u[27]^u[23]^u[21]^u[17]^u[16]^u[15]^u[12]^u[8]^u[7]^u[6]^u[5]^u[3]^u[0];
	y[241] = x[177]^x[236]^x[238]^x[240]^x[242]^x[243]^x[244]^x[245]^x[246]^x[249]^x[250]^x[256]^x[258]^x[260]^x[261]^x[264]^x[267]^x[269]^x[270]^x[271]^x[272]^x[273]^x[276]^x[277]^x[280]^x[283]^x[284]^x[287]^x[288]^x[289]^x[297]^x[298]^u[63]^u[61]^u[59]^u[57]^u[56]^u[55]^u[54]^u[53]^u[50]^u[49]^u[43]^u[41]^u[39]^u[38]^u[35]^u[32]^u[30]^u[29]^u[28]^u[27]^u[26]^u[23]^u[22]^u[19]^u[16]^u[15]^u[12]^u[11]^u[10]^u[2]^u[1];
	y[242] = x[178]^x[237]^x[239]^x[241]^x[243]^x[244]^x[245]^x[246]^x[247]^x[250]^x[251]^x[257]^x[259]^x[261]^x[262]^x[265]^x[268]^x[270]^x[271]^x[272]^x[273]^x[274]^x[277]^x[278]^x[281]^x[284]^x[285]^x[288]^x[289]^x[290]^x[298]^x[299]^u[62]^u[60]^u[58]^u[56]^u[55]^u[54]^u[53]^u[52]^u[49]^u[48]^u[42]^u[40]^u[38]^u[37]^u[34]^u[31]^u[29]^u[28]^u[27]^u[26]^u[25]^u[22]^u[21]^u[18]^u[15]^u[14]^u[11]^u[10]^u[9]^u[1]^u[0];
	y[243] = x[179]^x[238]^x[240]^x[242]^x[244]^x[245]^x[246]^x[247]^x[248]^x[251]^x[252]^x[258]^x[260]^x[262]^x[263]^x[266]^x[269]^x[271]^x[272]^x[273]^x[274]^x[275]^x[278]^x[279]^x[282]^x[285]^x[286]^x[289]^x[290]^x[291]^x[299]^u[61]^u[59]^u[57]^u[55]^u[54]^u[53]^u[52]^u[51]^u[48]^u[47]^u[41]^u[39]^u[37]^u[36]^u[33]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[21]^u[20]^u[17]^u[14]^u[13]^u[10]^u[9]^u[8]^u[0];
	y[244] = x[180]^x[239]^x[241]^x[243]^x[245]^x[246]^x[247]^x[248]^x[249]^x[252]^x[253]^x[259]^x[261]^x[263]^x[264]^x[267]^x[270]^x[272]^x[273]^x[274]^x[275]^x[276]^x[279]^x[280]^x[283]^x[286]^x[287]^x[290]^x[291]^x[292]^u[60]^u[58]^u[56]^u[54]^u[53]^u[52]^u[51]^u[50]^u[47]^u[46]^u[40]^u[38]^u[36]^u[35]^u[32]^u[29]^u[27]^u[26]^u[25]^u[24]^u[23]^u[20]^u[19]^u[16]^u[13]^u[12]^u[9]^u[8]^u[7];
	y[245] = x[181]^x[236]^x[238]^x[239]^x[240]^x[241]^x[242]^x[244]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[253]^x[254]^x[255]^x[262]^x[265]^x[268]^x[269]^x[273]^x[274]^x[275]^x[277]^x[279]^x[281]^x[284]^x[285]^x[288]^x[289]^x[291]^x[294]^x[295]^x[298]^u[63]^u[61]^u[60]^u[59]^u[58]^u[57]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[46]^u[45]^u[44]^u[37]^u[34]^u[31]^u[30]^u[26]^u[25]^u[24]^u[22]^u[20]^u[18]^u[15]^u[14]^u[11]^u[10]^u[8]^u[5]^u[4]^u[1];
	y[246] = x[182]^x[237]^x[239]^x[240]^x[241]^x[242]^x[243]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[254]^x[255]^x[256]^x[263]^x[266]^x[269]^x[270]^x[274]^x[275]^x[276]^x[278]^x[280]^x[282]^x[285]^x[286]^x[289]^x[290]^x[292]^x[295]^x[296]^x[299]^u[62]^u[60]^u[59]^u[58]^u[57]^u[56]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[45]^u[44]^u[43]^u[36]^u[33]^u[30]^u[29]^u[25]^u[24]^u[23]^u[21]^u[19]^u[17]^u[14]^u[13]^u[10]^u[9]^u[7]^u[4]^u[3]^u[0];
	y[247] = x[183]^x[236]^x[239]^x[240]^x[242]^x[243]^x[244]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[256]^x[257]^x[260]^x[267]^x[269]^x[270]^x[275]^x[277]^x[280]^x[281]^x[283]^x[285]^x[286]^x[289]^x[290]^x[291]^x[292]^x[294]^x[295]^x[296]^x[297]^x[298]^u[63]^u[60]^u[59]^u[57]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[43]^u[42]^u[39]^u[32]^u[30]^u[29]^u[24]^u[22]^u[19]^u[18]^u[16]^u[14]^u[13]^u[10]^u[9]^u[8]^u[7]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[248] = x[184]^x[237]^x[240]^x[241]^x[243]^x[244]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[257]^x[258]^x[261]^x[268]^x[270]^x[271]^x[276]^x[278]^x[281]^x[282]^x[284]^x[286]^x[287]^x[290]^x[291]^x[292]^x[293]^x[295]^x[296]^x[297]^x[298]^x[299]^u[62]^u[59]^u[58]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[42]^u[41]^u[38]^u[31]^u[29]^u[28]^u[23]^u[21]^u[18]^u[17]^u[15]^u[13]^u[12]^u[9]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[249] = x[185]^x[238]^x[241]^x[242]^x[244]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[258]^x[259]^x[262]^x[269]^x[271]^x[272]^x[277]^x[279]^x[282]^x[283]^x[285]^x[287]^x[288]^x[291]^x[292]^x[293]^x[294]^x[296]^x[297]^x[298]^x[299]^u[61]^u[58]^u[57]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[41]^u[40]^u[37]^u[30]^u[28]^u[27]^u[22]^u[20]^u[17]^u[16]^u[14]^u[12]^u[11]^u[8]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[250] = x[186]^x[239]^x[242]^x[243]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[255]^x[259]^x[260]^x[263]^x[270]^x[272]^x[273]^x[278]^x[280]^x[283]^x[284]^x[286]^x[288]^x[289]^x[292]^x[293]^x[294]^x[295]^x[297]^x[298]^x[299]^u[60]^u[57]^u[56]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[44]^u[40]^u[39]^u[36]^u[29]^u[27]^u[26]^u[21]^u[19]^u[16]^u[15]^u[13]^u[11]^u[10]^u[7]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[251] = x[187]^x[236]^x[238]^x[239]^x[240]^x[241]^x[243]^x[244]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[256]^x[261]^x[269]^x[273]^x[274]^x[276]^x[280]^x[281]^x[284]^x[290]^x[292]^x[296]^x[299]^u[63]^u[61]^u[60]^u[59]^u[58]^u[56]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[43]^u[38]^u[30]^u[26]^u[25]^u[23]^u[19]^u[18]^u[15]^u[9]^u[7]^u[3]^u[0];
	y[252] = x[188]^x[237]^x[239]^x[240]^x[241]^x[242]^x[244]^x[245]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[255]^x[257]^x[262]^x[270]^x[274]^x[275]^x[277]^x[281]^x[282]^x[285]^x[291]^x[293]^x[297]^u[62]^u[60]^u[59]^u[58]^u[57]^u[55]^u[54]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[44]^u[42]^u[37]^u[29]^u[25]^u[24]^u[22]^u[18]^u[17]^u[14]^u[8]^u[6]^u[2];
	y[253] = x[189]^x[236]^x[239]^x[240]^x[242]^x[243]^x[246]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[256]^x[258]^x[260]^x[263]^x[264]^x[269]^x[275]^x[278]^x[279]^x[280]^x[282]^x[283]^x[285]^x[286]^x[287]^x[289]^x[293]^x[295]^u[63]^u[60]^u[59]^u[57]^u[56]^u[53]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[43]^u[41]^u[39]^u[36]^u[35]^u[30]^u[24]^u[21]^u[20]^u[19]^u[17]^u[16]^u[14]^u[13]^u[12]^u[10]^u[6]^u[4];
	y[254] = x[190]^x[236]^x[237]^x[238]^x[239]^x[240]^x[243]^x[244]^x[245]^x[247]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[257]^x[259]^x[260]^x[261]^x[265]^x[269]^x[270]^x[271]^x[281]^x[283]^x[284]^x[285]^x[286]^x[288]^x[289]^x[290]^x[292]^x[293]^x[295]^x[296]^x[298]^u[63]^u[62]^u[61]^u[60]^u[59]^u[56]^u[55]^u[54]^u[52]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[42]^u[40]^u[39]^u[38]^u[34]^u[30]^u[29]^u[28]^u[18]^u[16]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[7]^u[6]^u[4]^u[3]^u[1];
	y[255] = x[191]^x[236]^x[237]^x[240]^x[244]^x[246]^x[248]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[258]^x[261]^x[262]^x[264]^x[266]^x[269]^x[270]^x[272]^x[276]^x[279]^x[280]^x[282]^x[284]^x[286]^x[290]^x[291]^x[292]^x[295]^x[296]^x[297]^x[298]^x[299]^u[63]^u[62]^u[59]^u[55]^u[53]^u[51]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[41]^u[38]^u[37]^u[35]^u[33]^u[30]^u[29]^u[27]^u[23]^u[20]^u[19]^u[17]^u[15]^u[13]^u[9]^u[8]^u[7]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[256] = x[192]^x[236]^x[237]^x[239]^x[247]^x[249]^x[250]^x[251]^x[252]^x[253]^x[254]^x[259]^x[260]^x[262]^x[263]^x[264]^x[265]^x[267]^x[269]^x[270]^x[273]^x[276]^x[277]^x[279]^x[281]^x[283]^x[289]^x[291]^x[294]^x[295]^x[296]^x[297]^x[299]^u[63]^u[62]^u[60]^u[52]^u[50]^u[49]^u[48]^u[47]^u[46]^u[45]^u[40]^u[39]^u[37]^u[36]^u[35]^u[34]^u[32]^u[30]^u[29]^u[26]^u[23]^u[22]^u[20]^u[18]^u[16]^u[10]^u[8]^u[5]^u[4]^u[3]^u[2]^u[0];
	y[257] = x[193]^x[237]^x[238]^x[240]^x[248]^x[250]^x[251]^x[252]^x[253]^x[254]^x[255]^x[260]^x[261]^x[263]^x[264]^x[265]^x[266]^x[268]^x[270]^x[271]^x[274]^x[277]^x[278]^x[280]^x[282]^x[284]^x[290]^x[292]^x[295]^x[296]^x[297]^x[298]^u[62]^u[61]^u[59]^u[51]^u[49]^u[48]^u[47]^u[46]^u[45]^u[44]^u[39]^u[38]^u[36]^u[35]^u[34]^u[33]^u[31]^u[29]^u[28]^u[25]^u[22]^u[21]^u[19]^u[17]^u[15]^u[9]^u[7]^u[4]^u[3]^u[2]^u[1];
	y[258] = x[194]^x[238]^x[239]^x[241]^x[249]^x[251]^x[252]^x[253]^x[254]^x[255]^x[256]^x[261]^x[262]^x[264]^x[265]^x[266]^x[267]^x[269]^x[271]^x[272]^x[275]^x[278]^x[279]^x[281]^x[283]^x[285]^x[291]^x[293]^x[296]^x[297]^x[298]^x[299]^u[61]^u[60]^u[58]^u[50]^u[48]^u[47]^u[46]^u[45]^u[44]^u[43]^u[38]^u[37]^u[35]^u[34]^u[33]^u[32]^u[30]^u[28]^u[27]^u[24]^u[21]^u[20]^u[18]^u[16]^u[14]^u[8]^u[6]^u[3]^u[2]^u[1]^u[0];
	y[259] = x[195]^x[236]^x[238]^x[240]^x[241]^x[242]^x[245]^x[250]^x[252]^x[253]^x[254]^x[256]^x[257]^x[260]^x[262]^x[263]^x[264]^x[265]^x[266]^x[267]^x[268]^x[269]^x[270]^x[271]^x[272]^x[273]^x[282]^x[284]^x[285]^x[286]^x[287]^x[289]^x[293]^x[295]^x[297]^x[299]^u[63]^u[61]^u[59]^u[58]^u[57]^u[54]^u[49]^u[47]^u[46]^u[45]^u[43]^u[42]^u[39]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[17]^u[15]^u[14]^u[13]^u[12]^u[10]^u[6]^u[4]^u[2]^u[0];
	y[260] = x[196]^x[236]^x[237]^x[238]^x[242]^x[243]^x[245]^x[246]^x[251]^x[253]^x[254]^x[257]^x[258]^x[260]^x[261]^x[263]^x[265]^x[266]^x[267]^x[268]^x[270]^x[272]^x[273]^x[274]^x[276]^x[279]^x[280]^x[283]^x[286]^x[288]^x[289]^x[290]^x[292]^x[293]^x[295]^x[296]^u[63]^u[62]^u[61]^u[57]^u[56]^u[54]^u[53]^u[48]^u[46]^u[45]^u[42]^u[41]^u[39]^u[38]^u[36]^u[34]^u[33]^u[32]^u[31]^u[29]^u[27]^u[26]^u[25]^u[23]^u[20]^u[19]^u[16]^u[13]^u[11]^u[10]^u[9]^u[7]^u[6]^u[4]^u[3];
	y[261] = x[197]^x[236]^x[237]^x[241]^x[243]^x[244]^x[245]^x[246]^x[247]^x[252]^x[254]^x[258]^x[259]^x[260]^x[261]^x[262]^x[266]^x[267]^x[268]^x[273]^x[274]^x[275]^x[276]^x[277]^x[279]^x[281]^x[284]^x[285]^x[290]^x[291]^x[292]^x[295]^x[296]^x[297]^x[298]^u[63]^u[62]^u[58]^u[56]^u[55]^u[54]^u[53]^u[52]^u[47]^u[45]^u[41]^u[40]^u[39]^u[38]^u[37]^u[33]^u[32]^u[31]^u[26]^u[25]^u[24]^u[23]^u[22]^u[20]^u[18]^u[15]^u[14]^u[9]^u[8]^u[7]^u[4]^u[3]^u[2]^u[1];
	y[262] = x[198]^x[237]^x[238]^x[242]^x[244]^x[245]^x[246]^x[247]^x[248]^x[253]^x[255]^x[259]^x[260]^x[261]^x[262]^x[263]^x[267]^x[268]^x[269]^x[274]^x[275]^x[276]^x[277]^x[278]^x[280]^x[282]^x[285]^x[286]^x[291]^x[292]^x[293]^x[296]^x[297]^x[298]^x[299]^u[62]^u[61]^u[57]^u[55]^u[54]^u[53]^u[52]^u[51]^u[46]^u[44]^u[40]^u[39]^u[38]^u[37]^u[36]^u[32]^u[31]^u[30]^u[25]^u[24]^u[23]^u[22]^u[21]^u[19]^u[17]^u[14]^u[13]^u[8]^u[7]^u[6]^u[3]^u[2]^u[1]^u[0];
	y[263] = x[199]^x[238]^x[239]^x[243]^x[245]^x[246]^x[247]^x[248]^x[249]^x[254]^x[256]^x[260]^x[261]^x[262]^x[263]^x[264]^x[268]^x[269]^x[270]^x[275]^x[276]^x[277]^x[278]^x[279]^x[281]^x[283]^x[286]^x[287]^x[292]^x[293]^x[294]^x[297]^x[298]^x[299]^u[61]^u[60]^u[56]^u[54]^u[53]^u[52]^u[51]^u[50]^u[45]^u[43]^u[39]^u[38]^u[37]^u[36]^u[35]^u[31]^u[30]^u[29]^u[24]^u[23]^u[22]^u[21]^u[20]^u[18]^u[16]^u[13]^u[12]^u[7]^u[6]^u[5]^u[2]^u[1]^u[0];
	y[264] = x[200]^x[239]^x[240]^x[244]^x[246]^x[247]^x[248]^x[249]^x[250]^x[255]^x[257]^x[261]^x[262]^x[263]^x[264]^x[265]^x[269]^x[270]^x[271]^x[276]^x[277]^x[278]^x[279]^x[280]^x[282]^x[284]^x[287]^x[288]^x[293]^x[294]^x[295]^x[298]^x[299]^u[60]^u[59]^u[55]^u[53]^u[52]^u[51]^u[50]^u[49]^u[44]^u[42]^u[38]^u[37]^u[36]^u[35]^u[34]^u[30]^u[29]^u[28]^u[23]^u[22]^u[21]^u[20]^u[19]^u[17]^u[15]^u[12]^u[11]^u[6]^u[5]^u[4]^u[1]^u[0];
	y[265] = x[201]^x[236]^x[238]^x[239]^x[240]^x[247]^x[248]^x[249]^x[250]^x[251]^x[255]^x[256]^x[258]^x[260]^x[262]^x[263]^x[265]^x[266]^x[269]^x[270]^x[272]^x[276]^x[277]^x[278]^x[281]^x[283]^x[287]^x[288]^x[292]^x[293]^x[296]^x[298]^x[299]^u[63]^u[61]^u[60]^u[59]^u[52]^u[51]^u[50]^u[49]^u[48]^u[44]^u[43]^u[41]^u[39]^u[37]^u[36]^u[34]^u[33]^u[30]^u[29]^u[27]^u[23]^u[22]^u[21]^u[18]^u[16]^u[12]^u[11]^u[7]^u[6]^u[3]^u[1]^u[0];
	y[266] = x[202]^x[236]^x[237]^x[238]^x[240]^x[245]^x[248]^x[249]^x[250]^x[251]^x[252]^x[255]^x[256]^x[257]^x[259]^x[260]^x[261]^x[263]^x[266]^x[267]^x[269]^x[270]^x[273]^x[276]^x[277]^x[278]^x[280]^x[282]^x[284]^x[285]^x[287]^x[288]^x[292]^x[295]^x[297]^x[298]^x[299]^u[63]^u[62]^u[61]^u[59]^u[54]^u[51]^u[50]^u[49]^u[48]^u[47]^u[44]^u[43]^u[42]^u[40]^u[39]^u[38]^u[36]^u[33]^u[32]^u[30]^u[29]^u[26]^u[23]^u[22]^u[21]^u[19]^u[17]^u[15]^u[14]^u[12]^u[11]^u[7]^u[4]^u[2]^u[1]^u[0];
	y[267] = x[203]^x[237]^x[238]^x[239]^x[241]^x[246]^x[249]^x[250]^x[251]^x[252]^x[253]^x[256]^x[257]^x[258]^x[260]^x[261]^x[262]^x[264]^x[267]^x[268]^x[270]^x[271]^x[274]^x[277]^x[278]^x[279]^x[281]^x[283]^x[285]^x[286]^x[288]^x[289]^x[293]^x[296]^x[298]^x[299]^u[62]^u[61]^u[60]^u[58]^u[53]^u[50]^u[49]^u[48]^u[47]^u[46]^u[43]^u[42]^u[41]^u[39]^u[38]^u[37]^u[35]^u[32]^u[31]^u[29]^u[28]^u[25]^u[22]^u[21]^u[20]^u[18]^u[16]^u[14]^u[13]^u[11]^u[10]^u[6]^u[3]^u[1]^u[0];
	y[268] = x[204]^x[236]^x[240]^x[241]^x[242]^x[245]^x[247]^x[250]^x[251]^x[252]^x[253]^x[254]^x[255]^x[257]^x[258]^x[259]^x[260]^x[261]^x[262]^x[263]^x[264]^x[265]^x[268]^x[272]^x[275]^x[276]^x[278]^x[282]^x[284]^x[285]^x[286]^x[290]^x[292]^x[293]^x[295]^x[297]^x[298]^x[299]^u[63]^u[59]^u[58]^u[57]^u[54]^u[52]^u[49]^u[48]^u[47]^u[46]^u[45]^u[44]^u[42]^u[41]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[31]^u[27]^u[24]^u[23]^u[21]^u[17]^u[15]^u[14]^u[13]^u[9]^u[7]^u[6]^u[4]^u[2]^u[1]^u[0];
	y[269] = x[205]^x[237]^x[241]^x[242]^x[243]^x[246]^x[248]^x[251]^x[252]^x[253]^x[254]^x[255]^x[256]^x[258]^x[259]^x[260]^x[261]^x[262]^x[263]^x[264]^x[265]^x[266]^x[269]^x[273]^x[276]^x[277]^x[279]^x[283]^x[285]^x[286]^x[287]^x[291]^x[293]^x[294]^x[296]^x[298]^x[299]^u[62]^u[58]^u[57]^u[56]^u[53]^u[51]^u[48]^u[47]^u[46]^u[45]^u[44]^u[43]^u[41]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[30]^u[26]^u[23]^u[22]^u[20]^u[16]^u[14]^u[13]^u[12]^u[8]^u[6]^u[5]^u[3]^u[1]^u[0];
	y[270] = x[206]^x[238]^x[242]^x[243]^x[244]^x[247]^x[249]^x[252]^x[253]^x[254]^x[255]^x[256]^x[257]^x[259]^x[260]^x[261]^x[262]^x[263]^x[264]^x[265]^x[266]^x[267]^x[270]^x[274]^x[277]^x[278]^x[280]^x[284]^x[286]^x[287]^x[288]^x[292]^x[294]^x[295]^x[297]^x[299]^u[61]^u[57]^u[56]^u[55]^u[52]^u[50]^u[47]^u[46]^u[45]^u[44]^u[43]^u[42]^u[40]^u[39]^u[38]^u[37]^u[36]^u[35]^u[34]^u[33]^u[32]^u[29]^u[25]^u[22]^u[21]^u[19]^u[15]^u[13]^u[12]^u[11]^u[7]^u[5]^u[4]^u[2]^u[0];
	y[271] = x[207]^x[236]^x[238]^x[241]^x[243]^x[244]^x[248]^x[250]^x[253]^x[254]^x[256]^x[257]^x[258]^x[261]^x[262]^x[263]^x[265]^x[266]^x[267]^x[268]^x[269]^x[275]^x[276]^x[278]^x[280]^x[281]^x[288]^x[292]^x[294]^x[296]^u[63]^u[61]^u[58]^u[56]^u[55]^u[51]^u[49]^u[46]^u[45]^u[43]^u[42]^u[41]^u[38]^u[37]^u[36]^u[34]^u[33]^u[32]^u[31]^u[30]^u[24]^u[23]^u[21]^u[19]^u[18]^u[11]^u[7]^u[5]^u[3];
	y[272] = x[208]^x[237]^x[239]^x[242]^x[244]^x[245]^x[249]^x[251]^x[254]^x[255]^x[257]^x[258]^x[259]^x[262]^x[263]^x[264]^x[266]^x[267]^x[268]^x[269]^x[270]^x[276]^x[277]^x[279]^x[281]^x[282]^x[289]^x[293]^x[295]^x[297]^u[62]^u[60]^u[57]^u[55]^u[54]^u[50]^u[48]^u[45]^u[44]^u[42]^u[41]^u[40]^u[37]^u[36]^u[35]^u[33]^u[32]^u[31]^u[30]^u[29]^u[23]^u[22]^u[20]^u[18]^u[17]^u[10]^u[6]^u[4]^u[2];
	y[273] = x[209]^x[236]^x[239]^x[240]^x[241]^x[243]^x[246]^x[250]^x[252]^x[256]^x[258]^x[259]^x[263]^x[265]^x[267]^x[268]^x[270]^x[276]^x[277]^x[278]^x[279]^x[282]^x[283]^x[285]^x[287]^x[289]^x[290]^x[292]^x[293]^x[295]^x[296]^u[63]^u[60]^u[59]^u[58]^u[56]^u[53]^u[49]^u[47]^u[43]^u[41]^u[40]^u[36]^u[34]^u[32]^u[31]^u[29]^u[23]^u[22]^u[21]^u[20]^u[17]^u[16]^u[14]^u[12]^u[10]^u[9]^u[7]^u[6]^u[4]^u[3];
	y[274] = x[210]^x[237]^x[240]^x[241]^x[242]^x[244]^x[247]^x[251]^x[253]^x[257]^x[259]^x[260]^x[264]^x[266]^x[268]^x[269]^x[271]^x[277]^x[278]^x[279]^x[280]^x[283]^x[284]^x[286]^x[288]^x[290]^x[291]^x[293]^x[294]^x[296]^x[297]^u[62]^u[59]^u[58]^u[57]^u[55]^u[52]^u[48]^u[46]^u[42]^u[40]^u[39]^u[35]^u[33]^u[31]^u[30]^u[28]^u[22]^u[21]^u[20]^u[19]^u[16]^u[15]^u[13]^u[11]^u[9]^u[8]^u[6]^u[5]^u[3]^u[2];
	y[275] = x[211]^x[236]^x[239]^x[242]^x[243]^x[248]^x[252]^x[254]^x[255]^x[258]^x[261]^x[264]^x[265]^x[267]^x[270]^x[271]^x[272]^x[276]^x[278]^x[281]^x[284]^x[291]^x[293]^x[297]^u[63]^u[60]^u[57]^u[56]^u[51]^u[47]^u[45]^u[44]^u[41]^u[38]^u[35]^u[34]^u[32]^u[29]^u[28]^u[27]^u[23]^u[21]^u[18]^u[15]^u[8]^u[6]^u[2];
	y[276] = x[212]^x[237]^x[240]^x[243]^x[244]^x[249]^x[253]^x[255]^x[256]^x[259]^x[262]^x[265]^x[266]^x[268]^x[271]^x[272]^x[273]^x[277]^x[279]^x[282]^x[285]^x[292]^x[294]^x[298]^u[62]^u[59]^u[56]^u[55]^u[50]^u[46]^u[44]^u[43]^u[40]^u[37]^u[34]^u[33]^u[31]^u[28]^u[27]^u[26]^u[22]^u[20]^u[17]^u[14]^u[7]^u[5]^u[1];
	y[277] = x[213]^x[236]^x[239]^x[244]^x[250]^x[254]^x[255]^x[256]^x[257]^x[263]^x[264]^x[266]^x[267]^x[271]^x[272]^x[273]^x[274]^x[276]^x[278]^x[279]^x[283]^x[285]^x[286]^x[287]^x[289]^x[292]^x[294]^x[298]^x[299]^u[63]^u[60]^u[55]^u[49]^u[45]^u[44]^u[43]^u[42]^u[36]^u[35]^u[33]^u[32]^u[28]^u[27]^u[26]^u[25]^u[23]^u[21]^u[20]^u[16]^u[14]^u[13]^u[12]^u[10]^u[7]^u[5]^u[1]^u[0];
	y[278] = x[214]^x[237]^x[240]^x[245]^x[251]^x[255]^x[256]^x[257]^x[258]^x[264]^x[265]^x[267]^x[268]^x[272]^x[273]^x[274]^x[275]^x[277]^x[279]^x[280]^x[284]^x[286]^x[287]^x[288]^x[290]^x[293]^x[295]^x[299]^u[62]^u[59]^u[54]^u[48]^u[44]^u[43]^u[42]^u[41]^u[35]^u[34]^u[32]^u[31]^u[27]^u[26]^u[25]^u[24]^u[22]^u[20]^u[19]^u[15]^u[13]^u[12]^u[11]^u[9]^u[6]^u[4]^u[0];
	y[279] = x[215]^x[236]^x[239]^x[245]^x[246]^x[252]^x[255]^x[256]^x[257]^x[258]^x[259]^x[260]^x[264]^x[265]^x[266]^x[268]^x[271]^x[273]^x[274]^x[275]^x[278]^x[279]^x[281]^x[288]^x[291]^x[292]^x[293]^x[295]^x[296]^x[298]^u[63]^u[60]^u[54]^u[53]^u[47]^u[44]^u[43]^u[42]^u[41]^u[40]^u[39]^u[35]^u[34]^u[33]^u[31]^u[28]^u[26]^u[25]^u[24]^u[21]^u[20]^u[18]^u[11]^u[8]^u[7]^u[6]^u[4]^u[3]^u[1];
	y[280] = x[216]^x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[245]^x[246]^x[247]^x[253]^x[255]^x[256]^x[257]^x[258]^x[259]^x[261]^x[264]^x[265]^x[266]^x[267]^x[271]^x[272]^x[274]^x[275]^x[282]^x[285]^x[287]^x[295]^x[296]^x[297]^x[298]^x[299]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[54]^u[53]^u[52]^u[46]^u[44]^u[43]^u[42]^u[41]^u[40]^u[38]^u[35]^u[34]^u[33]^u[32]^u[28]^u[27]^u[25]^u[24]^u[17]^u[14]^u[12]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[281] = x[217]^x[236]^x[237]^x[240]^x[242]^x[245]^x[246]^x[247]^x[248]^x[254]^x[255]^x[256]^x[257]^x[258]^x[259]^x[262]^x[264]^x[265]^x[266]^x[267]^x[268]^x[269]^x[271]^x[272]^x[273]^x[275]^x[279]^x[280]^x[283]^x[285]^x[286]^x[287]^x[288]^x[289]^x[292]^x[293]^x[294]^x[295]^x[296]^x[297]^x[299]^u[63]^u[62]^u[59]^u[57]^u[54]^u[53]^u[52]^u[51]^u[45]^u[44]^u[43]^u[42]^u[41]^u[40]^u[37]^u[35]^u[34]^u[33]^u[32]^u[31]^u[30]^u[28]^u[27]^u[26]^u[24]^u[20]^u[19]^u[16]^u[14]^u[13]^u[12]^u[11]^u[10]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2]^u[0];
	y[282] = x[218]^x[236]^x[237]^x[239]^x[243]^x[245]^x[246]^x[247]^x[248]^x[249]^x[256]^x[257]^x[258]^x[259]^x[263]^x[264]^x[265]^x[266]^x[267]^x[268]^x[270]^x[271]^x[272]^x[273]^x[274]^x[279]^x[281]^x[284]^x[285]^x[286]^x[288]^x[290]^x[292]^x[296]^x[297]^u[63]^u[62]^u[60]^u[56]^u[54]^u[53]^u[52]^u[51]^u[50]^u[43]^u[42]^u[41]^u[40]^u[36]^u[35]^u[34]^u[33]^u[32]^u[31]^u[29]^u[28]^u[27]^u[26]^u[25]^u[20]^u[18]^u[15]^u[14]^u[13]^u[11]^u[9]^u[7]^u[3]^u[2];
	y[283] = x[219]^x[237]^x[238]^x[240]^x[244]^x[246]^x[247]^x[248]^x[249]^x[250]^x[257]^x[258]^x[259]^x[260]^x[264]^x[265]^x[266]^x[267]^x[268]^x[269]^x[271]^x[272]^x[273]^x[274]^x[275]^x[280]^x[282]^x[285]^x[286]^x[287]^x[289]^x[291]^x[293]^x[297]^x[298]^u[62]^u[61]^u[59]^u[55]^u[53]^u[52]^u[51]^u[50]^u[49]^u[42]^u[41]^u[40]^u[39]^u[35]^u[34]^u[33]^u[32]^u[31]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[19]^u[17]^u[14]^u[13]^u[12]^u[10]^u[8]^u[6]^u[2]^u[1];
	y[284] = x[220]^x[236]^x[247]^x[248]^x[249]^x[250]^x[251]^x[255]^x[258]^x[259]^x[261]^x[264]^x[265]^x[266]^x[267]^x[268]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[279]^x[280]^x[281]^x[283]^x[285]^x[286]^x[288]^x[289]^x[290]^x[293]^x[295]^x[299]^u[63]^u[52]^u[51]^u[50]^u[49]^u[48]^u[44]^u[41]^u[40]^u[38]^u[35]^u[34]^u[33]^u[32]^u[31]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[20]^u[19]^u[18]^u[16]^u[14]^u[13]^u[11]^u[10]^u[9]^u[6]^u[4]^u[0];
	y[285] = x[221]^x[237]^x[248]^x[249]^x[250]^x[251]^x[252]^x[256]^x[259]^x[260]^x[262]^x[265]^x[266]^x[267]^x[268]^x[269]^x[271]^x[272]^x[273]^x[274]^x[275]^x[276]^x[280]^x[281]^x[282]^x[284]^x[286]^x[287]^x[289]^x[290]^x[291]^x[294]^x[296]^u[62]^u[51]^u[50]^u[49]^u[48]^u[47]^u[43]^u[40]^u[39]^u[37]^u[34]^u[33]^u[32]^u[31]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[19]^u[18]^u[17]^u[15]^u[13]^u[12]^u[10]^u[9]^u[8]^u[5]^u[3];
	y[286] = x[222]^x[236]^x[239]^x[241]^x[245]^x[249]^x[250]^x[251]^x[252]^x[253]^x[255]^x[257]^x[261]^x[263]^x[264]^x[266]^x[267]^x[268]^x[270]^x[271]^x[272]^x[273]^x[274]^x[275]^x[277]^x[279]^x[280]^x[281]^x[282]^x[283]^x[288]^x[289]^x[290]^x[291]^x[293]^x[294]^x[297]^x[298]^u[63]^u[60]^u[58]^u[54]^u[50]^u[49]^u[48]^u[47]^u[46]^u[44]^u[42]^u[38]^u[36]^u[35]^u[33]^u[32]^u[31]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[22]^u[20]^u[19]^u[18]^u[17]^u[16]^u[11]^u[10]^u[9]^u[8]^u[6]^u[5]^u[2]^u[1];
	y[287] = x[223]^x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[242]^x[245]^x[246]^x[250]^x[251]^x[252]^x[253]^x[254]^x[255]^x[256]^x[258]^x[260]^x[262]^x[265]^x[267]^x[268]^x[272]^x[273]^x[274]^x[275]^x[278]^x[279]^x[281]^x[282]^x[283]^x[284]^x[285]^x[287]^x[290]^x[291]^x[293]^x[299]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[57]^u[54]^u[53]^u[49]^u[48]^u[47]^u[46]^u[45]^u[44]^u[43]^u[41]^u[39]^u[37]^u[34]^u[32]^u[31]^u[27]^u[26]^u[25]^u[24]^u[21]^u[20]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[9]^u[8]^u[6]^u[0];
	y[288] = x[224]^x[236]^x[237]^x[240]^x[242]^x[243]^x[245]^x[246]^x[247]^x[251]^x[252]^x[253]^x[254]^x[256]^x[257]^x[259]^x[260]^x[261]^x[263]^x[264]^x[266]^x[268]^x[271]^x[273]^x[274]^x[275]^x[282]^x[283]^x[284]^x[286]^x[287]^x[288]^x[289]^x[291]^x[293]^x[295]^x[298]^u[63]^u[62]^u[59]^u[57]^u[56]^u[54]^u[53]^u[52]^u[48]^u[47]^u[46]^u[45]^u[43]^u[42]^u[40]^u[39]^u[38]^u[36]^u[35]^u[33]^u[31]^u[28]^u[26]^u[25]^u[24]^u[17]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[8]^u[6]^u[4]^u[1];
	y[289] = x[225]^x[237]^x[238]^x[241]^x[243]^x[244]^x[246]^x[247]^x[248]^x[252]^x[253]^x[254]^x[255]^x[257]^x[258]^x[260]^x[261]^x[262]^x[264]^x[265]^x[267]^x[269]^x[272]^x[274]^x[275]^x[276]^x[283]^x[284]^x[285]^x[287]^x[288]^x[289]^x[290]^x[292]^x[294]^x[296]^x[299]^u[62]^u[61]^u[58]^u[56]^u[55]^u[53]^u[52]^u[51]^u[47]^u[46]^u[45]^u[44]^u[42]^u[41]^u[39]^u[38]^u[37]^u[35]^u[34]^u[32]^u[30]^u[27]^u[25]^u[24]^u[23]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[7]^u[5]^u[3]^u[0];
	y[290] = x[226]^x[238]^x[239]^x[242]^x[244]^x[245]^x[247]^x[248]^x[249]^x[253]^x[254]^x[255]^x[256]^x[258]^x[259]^x[261]^x[262]^x[263]^x[265]^x[266]^x[268]^x[270]^x[273]^x[275]^x[276]^x[277]^x[284]^x[285]^x[286]^x[288]^x[289]^x[290]^x[291]^x[293]^x[295]^x[297]^u[61]^u[60]^u[57]^u[55]^u[54]^u[52]^u[51]^u[50]^u[46]^u[45]^u[44]^u[43]^u[41]^u[40]^u[38]^u[37]^u[36]^u[34]^u[33]^u[31]^u[29]^u[26]^u[24]^u[23]^u[22]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[6]^u[4]^u[2];
	y[291] = x[227]^x[236]^x[238]^x[240]^x[241]^x[243]^x[246]^x[248]^x[249]^x[250]^x[254]^x[256]^x[257]^x[259]^x[262]^x[263]^x[266]^x[267]^x[274]^x[277]^x[278]^x[279]^x[280]^x[286]^x[290]^x[291]^x[293]^x[295]^x[296]^u[63]^u[61]^u[59]^u[58]^u[56]^u[53]^u[51]^u[50]^u[49]^u[45]^u[43]^u[42]^u[40]^u[37]^u[36]^u[33]^u[32]^u[25]^u[22]^u[21]^u[20]^u[19]^u[13]^u[9]^u[8]^u[6]^u[4]^u[3];
	y[292] = x[228]^x[237]^x[239]^x[241]^x[242]^x[244]^x[247]^x[249]^x[250]^x[251]^x[255]^x[257]^x[258]^x[260]^x[263]^x[264]^x[267]^x[268]^x[275]^x[278]^x[279]^x[280]^x[281]^x[287]^x[291]^x[292]^x[294]^x[296]^x[297]^u[62]^u[60]^u[58]^u[57]^u[55]^u[52]^u[50]^u[49]^u[48]^u[44]^u[42]^u[41]^u[39]^u[36]^u[35]^u[32]^u[31]^u[24]^u[21]^u[20]^u[19]^u[18]^u[12]^u[8]^u[7]^u[5]^u[3]^u[2];
	y[293] = x[229]^x[236]^x[239]^x[240]^x[241]^x[242]^x[243]^x[248]^x[250]^x[251]^x[252]^x[255]^x[256]^x[258]^x[259]^x[260]^x[261]^x[265]^x[268]^x[271]^x[281]^x[282]^x[285]^x[287]^x[288]^x[289]^x[294]^x[297]^u[63]^u[60]^u[59]^u[58]^u[57]^u[56]^u[51]^u[49]^u[48]^u[47]^u[44]^u[43]^u[41]^u[40]^u[39]^u[38]^u[34]^u[31]^u[28]^u[18]^u[17]^u[14]^u[12]^u[11]^u[10]^u[5]^u[2];
	y[294] = x[230]^x[237]^x[240]^x[241]^x[242]^x[243]^x[244]^x[249]^x[251]^x[252]^x[253]^x[256]^x[257]^x[259]^x[260]^x[261]^x[262]^x[266]^x[269]^x[272]^x[282]^x[283]^x[286]^x[288]^x[289]^x[290]^x[295]^x[298]^u[62]^u[59]^u[58]^u[57]^u[56]^u[55]^u[50]^u[48]^u[47]^u[46]^u[43]^u[42]^u[40]^u[39]^u[38]^u[37]^u[33]^u[30]^u[27]^u[17]^u[16]^u[13]^u[11]^u[10]^u[9]^u[4]^u[1];
	y[295] = x[231]^x[236]^x[239]^x[242]^x[243]^x[244]^x[250]^x[252]^x[253]^x[254]^x[255]^x[257]^x[258]^x[261]^x[262]^x[263]^x[264]^x[267]^x[269]^x[270]^x[271]^x[273]^x[276]^x[279]^x[280]^x[283]^x[284]^x[285]^x[290]^x[291]^x[292]^x[293]^x[294]^x[295]^x[296]^x[298]^x[299]^u[63]^u[60]^u[57]^u[56]^u[55]^u[49]^u[47]^u[46]^u[45]^u[44]^u[42]^u[41]^u[38]^u[37]^u[36]^u[35]^u[32]^u[30]^u[29]^u[28]^u[26]^u[23]^u[20]^u[19]^u[16]^u[15]^u[14]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3]^u[1]^u[0];
	y[296] = x[232]^x[236]^x[237]^x[238]^x[239]^x[240]^x[241]^x[243]^x[244]^x[251]^x[253]^x[254]^x[256]^x[258]^x[259]^x[260]^x[262]^x[263]^x[265]^x[268]^x[269]^x[270]^x[272]^x[274]^x[276]^x[277]^x[279]^x[281]^x[284]^x[286]^x[287]^x[289]^x[291]^x[296]^x[297]^x[298]^x[299]^u[63]^u[62]^u[61]^u[60]^u[59]^u[58]^u[56]^u[55]^u[48]^u[46]^u[45]^u[43]^u[41]^u[40]^u[39]^u[37]^u[36]^u[34]^u[31]^u[30]^u[29]^u[27]^u[25]^u[23]^u[22]^u[20]^u[18]^u[15]^u[13]^u[12]^u[10]^u[8]^u[3]^u[2]^u[1]^u[0];
	y[297] = x[233]^x[236]^x[237]^x[240]^x[242]^x[244]^x[252]^x[254]^x[257]^x[259]^x[261]^x[263]^x[266]^x[270]^x[273]^x[275]^x[276]^x[277]^x[278]^x[279]^x[282]^x[288]^x[289]^x[290]^x[293]^x[294]^x[295]^x[297]^x[299]^u[63]^u[62]^u[59]^u[57]^u[55]^u[47]^u[45]^u[42]^u[40]^u[38]^u[36]^u[33]^u[29]^u[26]^u[24]^u[23]^u[22]^u[21]^u[20]^u[17]^u[11]^u[10]^u[9]^u[6]^u[5]^u[4]^u[2]^u[0];
	y[298] = x[234]^x[236]^x[237]^x[239]^x[243]^x[253]^x[258]^x[262]^x[267]^x[269]^x[274]^x[277]^x[278]^x[283]^x[285]^x[287]^x[290]^x[291]^x[292]^x[293]^x[296]^u[63]^u[62]^u[60]^u[56]^u[46]^u[41]^u[37]^u[32]^u[30]^u[25]^u[22]^u[21]^u[16]^u[14]^u[12]^u[9]^u[8]^u[7]^u[6]^u[3];
	y[299] = x[235]^x[237]^x[238]^x[240]^x[244]^x[254]^x[259]^x[263]^x[268]^x[270]^x[275]^x[278]^x[279]^x[284]^x[286]^x[288]^x[291]^x[292]^x[293]^x[294]^x[297]^u[62]^u[61]^u[59]^u[55]^u[45]^u[40]^u[36]^u[31]^u[29]^u[24]^u[21]^u[20]^u[15]^u[13]^u[11]^u[8]^u[7]^u[6]^u[5]^u[2];
	return y;
endfunction
