package BCH_common;

typedef Bit#(270) ENCODED;
typedef Bit#(64) MESSAGE;
typedef 256 MAX_MSG_IN_CNT_VAL;
typedef 10 MSG_IN_CNT_BIT_WIDTH; //16384/32
typedef 5 PARITY_CNT;
typedef 270 PARITY_LEN;
typedef Bit#(15) GF_SYM;
typedef 18 T_BCH; // error correcting capability
typedef 36 DOUBLE_T_BCH;
typedef Vector#(36, GF_SYM) SYNDROME;
typedef Vector#(19, GF_SYM) POLYNOMIAL;
typedef Vector#(19, GF_SYM) POLYNOMIAL_CHIEN;
typedef Int#(6) POLY_IDX;

typedef Bit#(64) EST_ERR_VEC;
typedef 64 PARALLELISM;

import Vector::*;
function Bit#(15) gf_add(Bit#(15) a, Bit#(15) b);
	return a ^ b;
endfunction

function Bit#(15) gf_div_prim_poly(Bit#(29) a);
	Bit#(15) a_q;
	a_q[0] = a[0]^a[15];
	a_q[1] = a[1]^a[15]^a[16];
	a_q[2] = a[2]^a[16]^a[17];
	a_q[3] = a[3]^a[17]^a[18];
	a_q[4] = a[4]^a[18]^a[19];
	a_q[5] = a[5]^a[19]^a[20];
	a_q[6] = a[6]^a[20]^a[21];
	a_q[7] = a[7]^a[21]^a[22];
	a_q[8] = a[8]^a[22]^a[23];
	a_q[9] = a[9]^a[23]^a[24];
	a_q[10] = a[10]^a[24]^a[25];
	a_q[11] = a[11]^a[25]^a[26];
	a_q[12] = a[12]^a[26]^a[27];
	a_q[13] = a[13]^a[27]^a[28];
	a_q[14] = a[14]^a[28];
	return a_q;
endfunction

(* noinline *)
function Bit#(15) gf_mul(Bit#(15) a, Bit#(15) b);
	Bit#(29) c;
	c[0] = (a[0] & b[0]);
	c[1] = (a[0] & b[1])^(a[1] & b[0]);
	c[2] = (a[0] & b[2])^(a[1] & b[1])^(a[2] & b[0]);
	c[3] = (a[0] & b[3])^(a[1] & b[2])^(a[2] & b[1])^(a[3] & b[0]);
	c[4] = (a[0] & b[4])^(a[1] & b[3])^(a[2] & b[2])^(a[3] & b[1])^(a[4] & b[0]);
	c[5] = (a[0] & b[5])^(a[1] & b[4])^(a[2] & b[3])^(a[3] & b[2])^(a[4] & b[1])^(a[5] & b[0]);
	c[6] = (a[0] & b[6])^(a[1] & b[5])^(a[2] & b[4])^(a[3] & b[3])^(a[4] & b[2])^(a[5] & b[1])^(a[6] & b[0]);
	c[7] = (a[0] & b[7])^(a[1] & b[6])^(a[2] & b[5])^(a[3] & b[4])^(a[4] & b[3])^(a[5] & b[2])^(a[6] & b[1])^(a[7] & b[0]);
	c[8] = (a[0] & b[8])^(a[1] & b[7])^(a[2] & b[6])^(a[3] & b[5])^(a[4] & b[4])^(a[5] & b[3])^(a[6] & b[2])^(a[7] & b[1])^(a[8] & b[0]);
	c[9] = (a[0] & b[9])^(a[1] & b[8])^(a[2] & b[7])^(a[3] & b[6])^(a[4] & b[5])^(a[5] & b[4])^(a[6] & b[3])^(a[7] & b[2])^(a[8] & b[1])^(a[9] & b[0]);
	c[10] = (a[0] & b[10])^(a[1] & b[9])^(a[2] & b[8])^(a[3] & b[7])^(a[4] & b[6])^(a[5] & b[5])^(a[6] & b[4])^(a[7] & b[3])^(a[8] & b[2])^(a[9] & b[1])^(a[10] & b[0]);
	c[11] = (a[0] & b[11])^(a[1] & b[10])^(a[2] & b[9])^(a[3] & b[8])^(a[4] & b[7])^(a[5] & b[6])^(a[6] & b[5])^(a[7] & b[4])^(a[8] & b[3])^(a[9] & b[2])^(a[10] & b[1])^(a[11] & b[0]);
	c[12] = (a[0] & b[12])^(a[1] & b[11])^(a[2] & b[10])^(a[3] & b[9])^(a[4] & b[8])^(a[5] & b[7])^(a[6] & b[6])^(a[7] & b[5])^(a[8] & b[4])^(a[9] & b[3])^(a[10] & b[2])^(a[11] & b[1])^(a[12] & b[0]);
	c[13] = (a[0] & b[13])^(a[1] & b[12])^(a[2] & b[11])^(a[3] & b[10])^(a[4] & b[9])^(a[5] & b[8])^(a[6] & b[7])^(a[7] & b[6])^(a[8] & b[5])^(a[9] & b[4])^(a[10] & b[3])^(a[11] & b[2])^(a[12] & b[1])^(a[13] & b[0]);
	c[14] = (a[0] & b[14])^(a[1] & b[13])^(a[2] & b[12])^(a[3] & b[11])^(a[4] & b[10])^(a[5] & b[9])^(a[6] & b[8])^(a[7] & b[7])^(a[8] & b[6])^(a[9] & b[5])^(a[10] & b[4])^(a[11] & b[3])^(a[12] & b[2])^(a[13] & b[1])^(a[14] & b[0]);
	c[15] = (a[1] & b[14])^(a[2] & b[13])^(a[3] & b[12])^(a[4] & b[11])^(a[5] & b[10])^(a[6] & b[9])^(a[7] & b[8])^(a[8] & b[7])^(a[9] & b[6])^(a[10] & b[5])^(a[11] & b[4])^(a[12] & b[3])^(a[13] & b[2])^(a[14] & b[1]);
	c[16] = (a[2] & b[14])^(a[3] & b[13])^(a[4] & b[12])^(a[5] & b[11])^(a[6] & b[10])^(a[7] & b[9])^(a[8] & b[8])^(a[9] & b[7])^(a[10] & b[6])^(a[11] & b[5])^(a[12] & b[4])^(a[13] & b[3])^(a[14] & b[2]);
	c[17] = (a[3] & b[14])^(a[4] & b[13])^(a[5] & b[12])^(a[6] & b[11])^(a[7] & b[10])^(a[8] & b[9])^(a[9] & b[8])^(a[10] & b[7])^(a[11] & b[6])^(a[12] & b[5])^(a[13] & b[4])^(a[14] & b[3]);
	c[18] = (a[4] & b[14])^(a[5] & b[13])^(a[6] & b[12])^(a[7] & b[11])^(a[8] & b[10])^(a[9] & b[9])^(a[10] & b[8])^(a[11] & b[7])^(a[12] & b[6])^(a[13] & b[5])^(a[14] & b[4]);
	c[19] = (a[5] & b[14])^(a[6] & b[13])^(a[7] & b[12])^(a[8] & b[11])^(a[9] & b[10])^(a[10] & b[9])^(a[11] & b[8])^(a[12] & b[7])^(a[13] & b[6])^(a[14] & b[5]);
	c[20] = (a[6] & b[14])^(a[7] & b[13])^(a[8] & b[12])^(a[9] & b[11])^(a[10] & b[10])^(a[11] & b[9])^(a[12] & b[8])^(a[13] & b[7])^(a[14] & b[6]);
	c[21] = (a[7] & b[14])^(a[8] & b[13])^(a[9] & b[12])^(a[10] & b[11])^(a[11] & b[10])^(a[12] & b[9])^(a[13] & b[8])^(a[14] & b[7]);
	c[22] = (a[8] & b[14])^(a[9] & b[13])^(a[10] & b[12])^(a[11] & b[11])^(a[12] & b[10])^(a[13] & b[9])^(a[14] & b[8]);
	c[23] = (a[9] & b[14])^(a[10] & b[13])^(a[11] & b[12])^(a[12] & b[11])^(a[13] & b[10])^(a[14] & b[9]);
	c[24] = (a[10] & b[14])^(a[11] & b[13])^(a[12] & b[12])^(a[13] & b[11])^(a[14] & b[10]);
	c[25] = (a[11] & b[14])^(a[12] & b[13])^(a[13] & b[12])^(a[14] & b[11]);
	c[26] = (a[12] & b[14])^(a[13] & b[13])^(a[14] & b[12]);
	c[27] = (a[13] & b[14])^(a[14] & b[13]);
	c[28] = (a[14] & b[14]);
	return gf_div_prim_poly(c);
endfunction


(* noinline *)
function Vector#(64, Bit#(15)) elp_evaluated(Vector#(19, Bit#(15)) reg_buffer);
	Vector#(64, Bit#(15)) elp_eval;
	elp_eval[0]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000000010)^gf_mul(reg_buffer[2], 15'b000000000000100)^gf_mul(reg_buffer[3], 15'b000000000001000)^gf_mul(reg_buffer[4], 15'b000000000010000)^gf_mul(reg_buffer[5], 15'b000000000100000)^gf_mul(reg_buffer[6], 15'b000000001000000)^gf_mul(reg_buffer[7], 15'b000000010000000)^gf_mul(reg_buffer[8], 15'b000000100000000)^gf_mul(reg_buffer[9], 15'b000001000000000)^gf_mul(reg_buffer[10], 15'b000010000000000)^gf_mul(reg_buffer[11], 15'b000100000000000)^gf_mul(reg_buffer[12], 15'b001000000000000)^gf_mul(reg_buffer[13], 15'b010000000000000)^gf_mul(reg_buffer[14], 15'b100000000000000)^gf_mul(reg_buffer[15], 15'b000000000000011)^gf_mul(reg_buffer[16], 15'b000000000000110)^gf_mul(reg_buffer[17], 15'b000000000001100)^gf_mul(reg_buffer[18], 15'b000000000011000);
	elp_eval[1]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000000100)^gf_mul(reg_buffer[2], 15'b000000000010000)^gf_mul(reg_buffer[3], 15'b000000001000000)^gf_mul(reg_buffer[4], 15'b000000100000000)^gf_mul(reg_buffer[5], 15'b000010000000000)^gf_mul(reg_buffer[6], 15'b001000000000000)^gf_mul(reg_buffer[7], 15'b100000000000000)^gf_mul(reg_buffer[8], 15'b000000000000110)^gf_mul(reg_buffer[9], 15'b000000000011000)^gf_mul(reg_buffer[10], 15'b000000001100000)^gf_mul(reg_buffer[11], 15'b000000110000000)^gf_mul(reg_buffer[12], 15'b000011000000000)^gf_mul(reg_buffer[13], 15'b001100000000000)^gf_mul(reg_buffer[14], 15'b110000000000000)^gf_mul(reg_buffer[15], 15'b000000000000101)^gf_mul(reg_buffer[16], 15'b000000000010100)^gf_mul(reg_buffer[17], 15'b000000001010000)^gf_mul(reg_buffer[18], 15'b000000101000000);
	elp_eval[2]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000001000)^gf_mul(reg_buffer[2], 15'b000000001000000)^gf_mul(reg_buffer[3], 15'b000001000000000)^gf_mul(reg_buffer[4], 15'b001000000000000)^gf_mul(reg_buffer[5], 15'b000000000000011)^gf_mul(reg_buffer[6], 15'b000000000011000)^gf_mul(reg_buffer[7], 15'b000000011000000)^gf_mul(reg_buffer[8], 15'b000011000000000)^gf_mul(reg_buffer[9], 15'b011000000000000)^gf_mul(reg_buffer[10], 15'b000000000000101)^gf_mul(reg_buffer[11], 15'b000000000101000)^gf_mul(reg_buffer[12], 15'b000000101000000)^gf_mul(reg_buffer[13], 15'b000101000000000)^gf_mul(reg_buffer[14], 15'b101000000000000)^gf_mul(reg_buffer[15], 15'b000000000001111)^gf_mul(reg_buffer[16], 15'b000000001111000)^gf_mul(reg_buffer[17], 15'b000001111000000)^gf_mul(reg_buffer[18], 15'b001111000000000);
	elp_eval[3]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000010000)^gf_mul(reg_buffer[2], 15'b000000100000000)^gf_mul(reg_buffer[3], 15'b001000000000000)^gf_mul(reg_buffer[4], 15'b000000000000110)^gf_mul(reg_buffer[5], 15'b000000001100000)^gf_mul(reg_buffer[6], 15'b000011000000000)^gf_mul(reg_buffer[7], 15'b110000000000000)^gf_mul(reg_buffer[8], 15'b000000000010100)^gf_mul(reg_buffer[9], 15'b000000101000000)^gf_mul(reg_buffer[10], 15'b001010000000000)^gf_mul(reg_buffer[11], 15'b100000000000110)^gf_mul(reg_buffer[12], 15'b000000001111000)^gf_mul(reg_buffer[13], 15'b000011110000000)^gf_mul(reg_buffer[14], 15'b111100000000000)^gf_mul(reg_buffer[15], 15'b000000000010001)^gf_mul(reg_buffer[16], 15'b000000100010000)^gf_mul(reg_buffer[17], 15'b001000100000000)^gf_mul(reg_buffer[18], 15'b001000000000110);
	elp_eval[4]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000100000)^gf_mul(reg_buffer[2], 15'b000010000000000)^gf_mul(reg_buffer[3], 15'b000000000000011)^gf_mul(reg_buffer[4], 15'b000000001100000)^gf_mul(reg_buffer[5], 15'b000110000000000)^gf_mul(reg_buffer[6], 15'b000000000000101)^gf_mul(reg_buffer[7], 15'b000000010100000)^gf_mul(reg_buffer[8], 15'b001010000000000)^gf_mul(reg_buffer[9], 15'b000000000001111)^gf_mul(reg_buffer[10], 15'b000000111100000)^gf_mul(reg_buffer[11], 15'b011110000000000)^gf_mul(reg_buffer[12], 15'b000000000010001)^gf_mul(reg_buffer[13], 15'b000001000100000)^gf_mul(reg_buffer[14], 15'b100010000000000)^gf_mul(reg_buffer[15], 15'b000000000110011)^gf_mul(reg_buffer[16], 15'b000011001100000)^gf_mul(reg_buffer[17], 15'b100110000000011)^gf_mul(reg_buffer[18], 15'b000000001010101);
	elp_eval[5]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000001000000)^gf_mul(reg_buffer[2], 15'b001000000000000)^gf_mul(reg_buffer[3], 15'b000000000011000)^gf_mul(reg_buffer[4], 15'b000011000000000)^gf_mul(reg_buffer[5], 15'b000000000000101)^gf_mul(reg_buffer[6], 15'b000000101000000)^gf_mul(reg_buffer[7], 15'b101000000000000)^gf_mul(reg_buffer[8], 15'b000000001111000)^gf_mul(reg_buffer[9], 15'b001111000000000)^gf_mul(reg_buffer[10], 15'b000000000010001)^gf_mul(reg_buffer[11], 15'b000010001000000)^gf_mul(reg_buffer[12], 15'b001000000000110)^gf_mul(reg_buffer[13], 15'b000000110011000)^gf_mul(reg_buffer[14], 15'b110011000000000)^gf_mul(reg_buffer[15], 15'b000000001010101)^gf_mul(reg_buffer[16], 15'b001010101000000)^gf_mul(reg_buffer[17], 15'b101000000011110)^gf_mul(reg_buffer[18], 15'b000011111111000);
	elp_eval[6]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000010000000)^gf_mul(reg_buffer[2], 15'b100000000000000)^gf_mul(reg_buffer[3], 15'b000000011000000)^gf_mul(reg_buffer[4], 15'b110000000000000)^gf_mul(reg_buffer[5], 15'b000000010100000)^gf_mul(reg_buffer[6], 15'b101000000000000)^gf_mul(reg_buffer[7], 15'b000000011110000)^gf_mul(reg_buffer[8], 15'b111100000000000)^gf_mul(reg_buffer[9], 15'b000000010001000)^gf_mul(reg_buffer[10], 15'b100010000000000)^gf_mul(reg_buffer[11], 15'b000000011001100)^gf_mul(reg_buffer[12], 15'b110011000000000)^gf_mul(reg_buffer[13], 15'b000000010101010)^gf_mul(reg_buffer[14], 15'b101010100000000)^gf_mul(reg_buffer[15], 15'b000000011111111)^gf_mul(reg_buffer[16], 15'b111111110000000)^gf_mul(reg_buffer[17], 15'b100000010000001)^gf_mul(reg_buffer[18], 15'b100000001000000);
	elp_eval[7]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000100000000)^gf_mul(reg_buffer[2], 15'b000000000000110)^gf_mul(reg_buffer[3], 15'b000011000000000)^gf_mul(reg_buffer[4], 15'b000000000010100)^gf_mul(reg_buffer[5], 15'b001010000000000)^gf_mul(reg_buffer[6], 15'b000000001111000)^gf_mul(reg_buffer[7], 15'b111100000000000)^gf_mul(reg_buffer[8], 15'b000000100010000)^gf_mul(reg_buffer[9], 15'b001000000000110)^gf_mul(reg_buffer[10], 15'b000011001100000)^gf_mul(reg_buffer[11], 15'b110000000010100)^gf_mul(reg_buffer[12], 15'b001010101000000)^gf_mul(reg_buffer[13], 15'b100000001111110)^gf_mul(reg_buffer[14], 15'b111111110000000)^gf_mul(reg_buffer[15], 15'b000000100000001)^gf_mul(reg_buffer[16], 15'b000000100000110)^gf_mul(reg_buffer[17], 15'b000011000000110)^gf_mul(reg_buffer[18], 15'b000011000010100);
	elp_eval[8]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000001000000000)^gf_mul(reg_buffer[2], 15'b000000000011000)^gf_mul(reg_buffer[3], 15'b011000000000000)^gf_mul(reg_buffer[4], 15'b000000101000000)^gf_mul(reg_buffer[5], 15'b000000000001111)^gf_mul(reg_buffer[6], 15'b001111000000000)^gf_mul(reg_buffer[7], 15'b000000010001000)^gf_mul(reg_buffer[8], 15'b001000000000110)^gf_mul(reg_buffer[9], 15'b000110011000000)^gf_mul(reg_buffer[10], 15'b000000001010101)^gf_mul(reg_buffer[11], 15'b010101000000011)^gf_mul(reg_buffer[12], 15'b000011111111000)^gf_mul(reg_buffer[13], 15'b111000000100001)^gf_mul(reg_buffer[14], 15'b100000001000000)^gf_mul(reg_buffer[15], 15'b000001100000011)^gf_mul(reg_buffer[16], 15'b000011000010100)^gf_mul(reg_buffer[17], 15'b010100000101000)^gf_mul(reg_buffer[18], 15'b101000111100000);
	elp_eval[9]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000010000000000)^gf_mul(reg_buffer[2], 15'b000000001100000)^gf_mul(reg_buffer[3], 15'b000000000000101)^gf_mul(reg_buffer[4], 15'b001010000000000)^gf_mul(reg_buffer[5], 15'b000000111100000)^gf_mul(reg_buffer[6], 15'b000000000010001)^gf_mul(reg_buffer[7], 15'b100010000000000)^gf_mul(reg_buffer[8], 15'b000011001100000)^gf_mul(reg_buffer[9], 15'b000000001010101)^gf_mul(reg_buffer[10], 15'b101010000000110)^gf_mul(reg_buffer[11], 15'b001111111100000)^gf_mul(reg_buffer[12], 15'b000000100000001)^gf_mul(reg_buffer[13], 15'b000010000011000)^gf_mul(reg_buffer[14], 15'b110000001100000)^gf_mul(reg_buffer[15], 15'b000010100000101)^gf_mul(reg_buffer[16], 15'b001010001111000)^gf_mul(reg_buffer[17], 15'b110000111100101)^gf_mul(reg_buffer[18], 15'b001000100010001);
	elp_eval[10]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000100000000000)^gf_mul(reg_buffer[2], 15'b000000110000000)^gf_mul(reg_buffer[3], 15'b000000000101000)^gf_mul(reg_buffer[4], 15'b100000000000110)^gf_mul(reg_buffer[5], 15'b011110000000000)^gf_mul(reg_buffer[6], 15'b000010001000000)^gf_mul(reg_buffer[7], 15'b000000011001100)^gf_mul(reg_buffer[8], 15'b110000000010100)^gf_mul(reg_buffer[9], 15'b010101000000011)^gf_mul(reg_buffer[10], 15'b001111111100000)^gf_mul(reg_buffer[11], 15'b000001000000010)^gf_mul(reg_buffer[12], 15'b001000001100000)^gf_mul(reg_buffer[13], 15'b000001100001010)^gf_mul(reg_buffer[14], 15'b101000001010000)^gf_mul(reg_buffer[15], 15'b000111100001111)^gf_mul(reg_buffer[16], 15'b111100100010000)^gf_mul(reg_buffer[17], 15'b000100010110011)^gf_mul(reg_buffer[18], 15'b001100110011101);
	elp_eval[11]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b001000000000000)^gf_mul(reg_buffer[2], 15'b000011000000000)^gf_mul(reg_buffer[3], 15'b000000101000000)^gf_mul(reg_buffer[4], 15'b000000001111000)^gf_mul(reg_buffer[5], 15'b000000000010001)^gf_mul(reg_buffer[6], 15'b001000000000110)^gf_mul(reg_buffer[7], 15'b110011000000000)^gf_mul(reg_buffer[8], 15'b001010101000000)^gf_mul(reg_buffer[9], 15'b000011111111000)^gf_mul(reg_buffer[10], 15'b000000100000001)^gf_mul(reg_buffer[11], 15'b001000001100000)^gf_mul(reg_buffer[12], 15'b000011000010100)^gf_mul(reg_buffer[13], 15'b100000101000110)^gf_mul(reg_buffer[14], 15'b111100001111000)^gf_mul(reg_buffer[15], 15'b001000100010001)^gf_mul(reg_buffer[16], 15'b001011001100110)^gf_mul(reg_buffer[17], 15'b110011101010100)^gf_mul(reg_buffer[18], 15'b101010100111110);
	elp_eval[12]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b010000000000000)^gf_mul(reg_buffer[2], 15'b001100000000000)^gf_mul(reg_buffer[3], 15'b000101000000000)^gf_mul(reg_buffer[4], 15'b000011110000000)^gf_mul(reg_buffer[5], 15'b000001000100000)^gf_mul(reg_buffer[6], 15'b000000110011000)^gf_mul(reg_buffer[7], 15'b000000010101010)^gf_mul(reg_buffer[8], 15'b100000001111110)^gf_mul(reg_buffer[9], 15'b111000000100001)^gf_mul(reg_buffer[10], 15'b000010000011000)^gf_mul(reg_buffer[11], 15'b000001100001010)^gf_mul(reg_buffer[12], 15'b100000101000110)^gf_mul(reg_buffer[13], 15'b111000011110011)^gf_mul(reg_buffer[14], 15'b100010001000100)^gf_mul(reg_buffer[15], 15'b011001100110011)^gf_mul(reg_buffer[16], 15'b111010101010100)^gf_mul(reg_buffer[17], 15'b010011111111111)^gf_mul(reg_buffer[18], 15'b111101000000001);
	elp_eval[13]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b100000000000000)^gf_mul(reg_buffer[2], 15'b110000000000000)^gf_mul(reg_buffer[3], 15'b101000000000000)^gf_mul(reg_buffer[4], 15'b111100000000000)^gf_mul(reg_buffer[5], 15'b100010000000000)^gf_mul(reg_buffer[6], 15'b110011000000000)^gf_mul(reg_buffer[7], 15'b101010100000000)^gf_mul(reg_buffer[8], 15'b111111110000000)^gf_mul(reg_buffer[9], 15'b100000001000000)^gf_mul(reg_buffer[10], 15'b110000001100000)^gf_mul(reg_buffer[11], 15'b101000001010000)^gf_mul(reg_buffer[12], 15'b111100001111000)^gf_mul(reg_buffer[13], 15'b100010001000100)^gf_mul(reg_buffer[14], 15'b110011001100110)^gf_mul(reg_buffer[15], 15'b101010101010101)^gf_mul(reg_buffer[16], 15'b011111111111110)^gf_mul(reg_buffer[17], 15'b010000000000001)^gf_mul(reg_buffer[18], 15'b111000000000000);
	elp_eval[14]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000000011)^gf_mul(reg_buffer[2], 15'b000000000000101)^gf_mul(reg_buffer[3], 15'b000000000001111)^gf_mul(reg_buffer[4], 15'b000000000010001)^gf_mul(reg_buffer[5], 15'b000000000110011)^gf_mul(reg_buffer[6], 15'b000000001010101)^gf_mul(reg_buffer[7], 15'b000000011111111)^gf_mul(reg_buffer[8], 15'b000000100000001)^gf_mul(reg_buffer[9], 15'b000001100000011)^gf_mul(reg_buffer[10], 15'b000010100000101)^gf_mul(reg_buffer[11], 15'b000111100001111)^gf_mul(reg_buffer[12], 15'b001000100010001)^gf_mul(reg_buffer[13], 15'b011001100110011)^gf_mul(reg_buffer[14], 15'b101010101010101)^gf_mul(reg_buffer[15], 15'b111111111111100)^gf_mul(reg_buffer[16], 15'b000000000000111)^gf_mul(reg_buffer[17], 15'b000000000001001)^gf_mul(reg_buffer[18], 15'b000000000011011);
	elp_eval[15]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000000110)^gf_mul(reg_buffer[2], 15'b000000000010100)^gf_mul(reg_buffer[3], 15'b000000001111000)^gf_mul(reg_buffer[4], 15'b000000100010000)^gf_mul(reg_buffer[5], 15'b000011001100000)^gf_mul(reg_buffer[6], 15'b001010101000000)^gf_mul(reg_buffer[7], 15'b111111110000000)^gf_mul(reg_buffer[8], 15'b000000100000110)^gf_mul(reg_buffer[9], 15'b000011000010100)^gf_mul(reg_buffer[10], 15'b001010001111000)^gf_mul(reg_buffer[11], 15'b111100100010000)^gf_mul(reg_buffer[12], 15'b001011001100110)^gf_mul(reg_buffer[13], 15'b111010101010100)^gf_mul(reg_buffer[14], 15'b011111111111110)^gf_mul(reg_buffer[15], 15'b000000000000111)^gf_mul(reg_buffer[16], 15'b000000000010010)^gf_mul(reg_buffer[17], 15'b000000001101100)^gf_mul(reg_buffer[18], 15'b000000101101000);
	elp_eval[16]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000001100)^gf_mul(reg_buffer[2], 15'b000000001010000)^gf_mul(reg_buffer[3], 15'b000001111000000)^gf_mul(reg_buffer[4], 15'b001000100000000)^gf_mul(reg_buffer[5], 15'b100110000000011)^gf_mul(reg_buffer[6], 15'b101000000011110)^gf_mul(reg_buffer[7], 15'b100000010000001)^gf_mul(reg_buffer[8], 15'b000011000000110)^gf_mul(reg_buffer[9], 15'b010100000101000)^gf_mul(reg_buffer[10], 15'b110000111100101)^gf_mul(reg_buffer[11], 15'b000100010110011)^gf_mul(reg_buffer[12], 15'b110011101010100)^gf_mul(reg_buffer[13], 15'b010011111111111)^gf_mul(reg_buffer[14], 15'b010000000000001)^gf_mul(reg_buffer[15], 15'b000000000001001)^gf_mul(reg_buffer[16], 15'b000000001101100)^gf_mul(reg_buffer[17], 15'b000001011010000)^gf_mul(reg_buffer[18], 15'b001110111000000);
	elp_eval[17]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000011000)^gf_mul(reg_buffer[2], 15'b000000101000000)^gf_mul(reg_buffer[3], 15'b001111000000000)^gf_mul(reg_buffer[4], 15'b001000000000110)^gf_mul(reg_buffer[5], 15'b000000001010101)^gf_mul(reg_buffer[6], 15'b000011111111000)^gf_mul(reg_buffer[7], 15'b100000001000000)^gf_mul(reg_buffer[8], 15'b000011000010100)^gf_mul(reg_buffer[9], 15'b101000111100000)^gf_mul(reg_buffer[10], 15'b001000100010001)^gf_mul(reg_buffer[11], 15'b001100110011101)^gf_mul(reg_buffer[12], 15'b101010100111110)^gf_mul(reg_buffer[13], 15'b111101000000001)^gf_mul(reg_buffer[14], 15'b111000000000000)^gf_mul(reg_buffer[15], 15'b000000000011011)^gf_mul(reg_buffer[16], 15'b000000101101000)^gf_mul(reg_buffer[17], 15'b001110111000000)^gf_mul(reg_buffer[18], 15'b011001000000110);
	elp_eval[18]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000110000)^gf_mul(reg_buffer[2], 15'b000010100000000)^gf_mul(reg_buffer[3], 15'b111000000000011)^gf_mul(reg_buffer[4], 15'b000000001100110)^gf_mul(reg_buffer[5], 15'b000101010100000)^gf_mul(reg_buffer[6], 15'b111111000000101)^gf_mul(reg_buffer[7], 15'b010000011000000)^gf_mul(reg_buffer[8], 15'b001010000010100)^gf_mul(reg_buffer[9], 15'b100001111001001)^gf_mul(reg_buffer[10], 15'b100010110011000)^gf_mul(reg_buffer[11], 15'b110101010101011)^gf_mul(reg_buffer[12], 15'b111111111101001)^gf_mul(reg_buffer[13], 15'b000001110000000)^gf_mul(reg_buffer[14], 15'b100100000000000)^gf_mul(reg_buffer[15], 15'b000000000101101)^gf_mul(reg_buffer[16], 15'b000011101110000)^gf_mul(reg_buffer[17], 15'b001100100000011)^gf_mul(reg_buffer[18], 15'b011000001011111);
	elp_eval[19]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000001100000)^gf_mul(reg_buffer[2], 15'b001010000000000)^gf_mul(reg_buffer[3], 15'b000000000010001)^gf_mul(reg_buffer[4], 15'b000011001100000)^gf_mul(reg_buffer[5], 15'b101010000000110)^gf_mul(reg_buffer[6], 15'b000000100000001)^gf_mul(reg_buffer[7], 15'b110000001100000)^gf_mul(reg_buffer[8], 15'b001010001111000)^gf_mul(reg_buffer[9], 15'b001000100010001)^gf_mul(reg_buffer[10], 15'b110011001110100)^gf_mul(reg_buffer[11], 15'b101001111111110)^gf_mul(reg_buffer[12], 15'b000000000000111)^gf_mul(reg_buffer[13], 15'b000000100100000)^gf_mul(reg_buffer[14], 15'b110110000000000)^gf_mul(reg_buffer[15], 15'b000000001110111)^gf_mul(reg_buffer[16], 15'b001001100100000)^gf_mul(reg_buffer[17], 15'b010110000010111)^gf_mul(reg_buffer[18], 15'b000011100000111);
	elp_eval[20]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000011000000)^gf_mul(reg_buffer[2], 15'b101000000000000)^gf_mul(reg_buffer[3], 15'b000000010001000)^gf_mul(reg_buffer[4], 15'b110011000000000)^gf_mul(reg_buffer[5], 15'b000000011111111)^gf_mul(reg_buffer[6], 15'b100000001000000)^gf_mul(reg_buffer[7], 15'b011000010100000)^gf_mul(reg_buffer[8], 15'b111100001111000)^gf_mul(reg_buffer[9], 15'b010001011001100)^gf_mul(reg_buffer[10], 15'b101010101010101)^gf_mul(reg_buffer[11], 15'b111111101000001)^gf_mul(reg_buffer[12], 15'b111000000000000)^gf_mul(reg_buffer[13], 15'b000000011011000)^gf_mul(reg_buffer[14], 15'b101101000000000)^gf_mul(reg_buffer[15], 15'b000000010011001)^gf_mul(reg_buffer[16], 15'b110101011000000)^gf_mul(reg_buffer[17], 15'b101000011100001)^gf_mul(reg_buffer[18], 15'b100100001001000);
	elp_eval[21]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000110000000)^gf_mul(reg_buffer[2], 15'b100000000000110)^gf_mul(reg_buffer[3], 15'b000010001000000)^gf_mul(reg_buffer[4], 15'b110000000010100)^gf_mul(reg_buffer[5], 15'b001111111100000)^gf_mul(reg_buffer[6], 15'b001000001100000)^gf_mul(reg_buffer[7], 15'b101000001010000)^gf_mul(reg_buffer[8], 15'b111100100010000)^gf_mul(reg_buffer[9], 15'b001100110011101)^gf_mul(reg_buffer[10], 15'b101001111111110)^gf_mul(reg_buffer[11], 15'b000000000011100)^gf_mul(reg_buffer[12], 15'b001001000000000)^gf_mul(reg_buffer[13], 15'b000000001011010)^gf_mul(reg_buffer[14], 15'b111011100000000)^gf_mul(reg_buffer[15], 15'b000000110101011)^gf_mul(reg_buffer[16], 15'b111111010000110)^gf_mul(reg_buffer[17], 15'b100010010000101)^gf_mul(reg_buffer[18], 15'b100011011010111);
	elp_eval[22]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000001100000000)^gf_mul(reg_buffer[2], 15'b000000000011110)^gf_mul(reg_buffer[3], 15'b010001000000000)^gf_mul(reg_buffer[4], 15'b000000101010100)^gf_mul(reg_buffer[5], 15'b111110000001001)^gf_mul(reg_buffer[6], 15'b001100000011000)^gf_mul(reg_buffer[7], 15'b010100011110000)^gf_mul(reg_buffer[8], 15'b001000100010110)^gf_mul(reg_buffer[9], 15'b011101010101010)^gf_mul(reg_buffer[10], 15'b111111110100001)^gf_mul(reg_buffer[11], 15'b110000000000011)^gf_mul(reg_buffer[12], 15'b000011011000000)^gf_mul(reg_buffer[13], 15'b100000000111010)^gf_mul(reg_buffer[14], 15'b100110010000000)^gf_mul(reg_buffer[15], 15'b000001011111101)^gf_mul(reg_buffer[16], 15'b000011100010010)^gf_mul(reg_buffer[17], 15'b011011000110110)^gf_mul(reg_buffer[18], 15'b101101111011100);
	elp_eval[23]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000011000000000)^gf_mul(reg_buffer[2], 15'b000000001111000)^gf_mul(reg_buffer[3], 15'b001000000000110)^gf_mul(reg_buffer[4], 15'b001010101000000)^gf_mul(reg_buffer[5], 15'b000000100000001)^gf_mul(reg_buffer[6], 15'b000011000010100)^gf_mul(reg_buffer[7], 15'b111100001111000)^gf_mul(reg_buffer[8], 15'b001011001100110)^gf_mul(reg_buffer[9], 15'b101010100111110)^gf_mul(reg_buffer[10], 15'b000000000000111)^gf_mul(reg_buffer[11], 15'b001001000000000)^gf_mul(reg_buffer[12], 15'b000000101101000)^gf_mul(reg_buffer[13], 15'b111000000010010)^gf_mul(reg_buffer[14], 15'b110101011000000)^gf_mul(reg_buffer[15], 15'b000011100000111)^gf_mul(reg_buffer[16], 15'b001001001101100)^gf_mul(reg_buffer[17], 15'b110100101101110)^gf_mul(reg_buffer[18], 15'b110001100110010);
	elp_eval[24]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000110000000000)^gf_mul(reg_buffer[2], 15'b000000111100000)^gf_mul(reg_buffer[3], 15'b000000000110011)^gf_mul(reg_buffer[4], 15'b101010000000110)^gf_mul(reg_buffer[5], 15'b010000000100000)^gf_mul(reg_buffer[6], 15'b000010100000101)^gf_mul(reg_buffer[7], 15'b011110010001000)^gf_mul(reg_buffer[8], 15'b110011001110100)^gf_mul(reg_buffer[9], 15'b111111111111100)^gf_mul(reg_buffer[10], 15'b001110000000000)^gf_mul(reg_buffer[11], 15'b000001101100000)^gf_mul(reg_buffer[12], 15'b000000001110111)^gf_mul(reg_buffer[13], 15'b110010000001100)^gf_mul(reg_buffer[14], 15'b101111110100000)^gf_mul(reg_buffer[15], 15'b000100100001001)^gf_mul(reg_buffer[16], 15'b110110101101000)^gf_mul(reg_buffer[17], 15'b110111011000111)^gf_mul(reg_buffer[18], 15'b010101010101110);
	elp_eval[25]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b001100000000000)^gf_mul(reg_buffer[2], 15'b000011110000000)^gf_mul(reg_buffer[3], 15'b000000110011000)^gf_mul(reg_buffer[4], 15'b100000001111110)^gf_mul(reg_buffer[5], 15'b000010000011000)^gf_mul(reg_buffer[6], 15'b100000101000110)^gf_mul(reg_buffer[7], 15'b100010001000100)^gf_mul(reg_buffer[8], 15'b111010101010100)^gf_mul(reg_buffer[9], 15'b111101000000001)^gf_mul(reg_buffer[10], 15'b000000100100000)^gf_mul(reg_buffer[11], 15'b000000001011010)^gf_mul(reg_buffer[12], 15'b111000000010010)^gf_mul(reg_buffer[13], 15'b010101100000101)^gf_mul(reg_buffer[14], 15'b111000001110000)^gf_mul(reg_buffer[15], 15'b001101100011011)^gf_mul(reg_buffer[16], 15'b110111101110110)^gf_mul(reg_buffer[17], 15'b100110100101011)^gf_mul(reg_buffer[18], 15'b111111110011001);
	elp_eval[26]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b011000000000000)^gf_mul(reg_buffer[2], 15'b001111000000000)^gf_mul(reg_buffer[3], 15'b000110011000000)^gf_mul(reg_buffer[4], 15'b000011111111000)^gf_mul(reg_buffer[5], 15'b000001100000011)^gf_mul(reg_buffer[6], 15'b101000111100000)^gf_mul(reg_buffer[7], 15'b010001011001100)^gf_mul(reg_buffer[8], 15'b101010100111110)^gf_mul(reg_buffer[9], 15'b000000000111000)^gf_mul(reg_buffer[10], 15'b000000000011011)^gf_mul(reg_buffer[11], 15'b101000000001111)^gf_mul(reg_buffer[12], 15'b011001000000110)^gf_mul(reg_buffer[13], 15'b011111101000011)^gf_mul(reg_buffer[14], 15'b100100001001000)^gf_mul(reg_buffer[15], 15'b010110100101101)^gf_mul(reg_buffer[16], 15'b110001100110010)^gf_mul(reg_buffer[17], 15'b101110111111110)^gf_mul(reg_buffer[18], 15'b000010101000000);
	elp_eval[27]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b110000000000000)^gf_mul(reg_buffer[2], 15'b111100000000000)^gf_mul(reg_buffer[3], 15'b110011000000000)^gf_mul(reg_buffer[4], 15'b111111110000000)^gf_mul(reg_buffer[5], 15'b110000001100000)^gf_mul(reg_buffer[6], 15'b111100001111000)^gf_mul(reg_buffer[7], 15'b110011001100110)^gf_mul(reg_buffer[8], 15'b011111111111110)^gf_mul(reg_buffer[9], 15'b111000000000000)^gf_mul(reg_buffer[10], 15'b110110000000000)^gf_mul(reg_buffer[11], 15'b111011100000000)^gf_mul(reg_buffer[12], 15'b110101011000000)^gf_mul(reg_buffer[13], 15'b111000001110000)^gf_mul(reg_buffer[14], 15'b110110001101100)^gf_mul(reg_buffer[15], 15'b111011101110111)^gf_mul(reg_buffer[16], 15'b100101010101010)^gf_mul(reg_buffer[17], 15'b001100000000001)^gf_mul(reg_buffer[18], 15'b111111000000000);
	elp_eval[28]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b100000000000011)^gf_mul(reg_buffer[2], 15'b110000000000101)^gf_mul(reg_buffer[3], 15'b011000000001010)^gf_mul(reg_buffer[4], 15'b111100000010001)^gf_mul(reg_buffer[5], 15'b000110000101000)^gf_mul(reg_buffer[6], 15'b001111001000100)^gf_mul(reg_buffer[7], 15'b011001110101010)^gf_mul(reg_buffer[8], 15'b111111010000001)^gf_mul(reg_buffer[9], 15'b000001001000000)^gf_mul(reg_buffer[10], 15'b000010110100000)^gf_mul(reg_buffer[11], 15'b000100110010000)^gf_mul(reg_buffer[12], 15'b001011111101000)^gf_mul(reg_buffer[13], 15'b010010000100100)^gf_mul(reg_buffer[14], 15'b101101001011010)^gf_mul(reg_buffer[15], 15'b001100110011010)^gf_mul(reg_buffer[16], 15'b011111111111001)^gf_mul(reg_buffer[17], 15'b010000000001111)^gf_mul(reg_buffer[18], 15'b001000000011000);
	elp_eval[29]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000000101)^gf_mul(reg_buffer[2], 15'b000000000010001)^gf_mul(reg_buffer[3], 15'b000000001010101)^gf_mul(reg_buffer[4], 15'b000000100000001)^gf_mul(reg_buffer[5], 15'b000010100000101)^gf_mul(reg_buffer[6], 15'b001000100010001)^gf_mul(reg_buffer[7], 15'b101010101010101)^gf_mul(reg_buffer[8], 15'b000000000000111)^gf_mul(reg_buffer[9], 15'b000000000011011)^gf_mul(reg_buffer[10], 15'b000000001110111)^gf_mul(reg_buffer[11], 15'b000000110101011)^gf_mul(reg_buffer[12], 15'b000011100000111)^gf_mul(reg_buffer[13], 15'b001101100011011)^gf_mul(reg_buffer[14], 15'b111011101110111)^gf_mul(reg_buffer[15], 15'b010101010101110)^gf_mul(reg_buffer[16], 15'b000000000010101)^gf_mul(reg_buffer[17], 15'b000000001000001)^gf_mul(reg_buffer[18], 15'b000000101000101);
	elp_eval[30]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000001010)^gf_mul(reg_buffer[2], 15'b000000001000100)^gf_mul(reg_buffer[3], 15'b000001010101000)^gf_mul(reg_buffer[4], 15'b001000000010000)^gf_mul(reg_buffer[5], 15'b010000010100011)^gf_mul(reg_buffer[6], 15'b100010001011000)^gf_mul(reg_buffer[7], 15'b010101001111111)^gf_mul(reg_buffer[8], 15'b000011100000000)^gf_mul(reg_buffer[9], 15'b011011000000000)^gf_mul(reg_buffer[10], 15'b101110000000101)^gf_mul(reg_buffer[11], 15'b101100000101110)^gf_mul(reg_buffer[12], 15'b111000100100000)^gf_mul(reg_buffer[13], 15'b110101101001010)^gf_mul(reg_buffer[14], 15'b000110011001101)^gf_mul(reg_buffer[15], 15'b111111111110010)^gf_mul(reg_buffer[16], 15'b000000001111110)^gf_mul(reg_buffer[17], 15'b000001100001100)^gf_mul(reg_buffer[18], 15'b001111001111000);
	elp_eval[31]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000010100)^gf_mul(reg_buffer[2], 15'b000000100010000)^gf_mul(reg_buffer[3], 15'b001010101000000)^gf_mul(reg_buffer[4], 15'b000000100000110)^gf_mul(reg_buffer[5], 15'b001010001111000)^gf_mul(reg_buffer[6], 15'b001011001100110)^gf_mul(reg_buffer[7], 15'b011111111111110)^gf_mul(reg_buffer[8], 15'b000000000010010)^gf_mul(reg_buffer[9], 15'b000000101101000)^gf_mul(reg_buffer[10], 15'b001001100100000)^gf_mul(reg_buffer[11], 15'b111111010000110)^gf_mul(reg_buffer[12], 15'b001001001101100)^gf_mul(reg_buffer[13], 15'b110111101110110)^gf_mul(reg_buffer[14], 15'b100101010101010)^gf_mul(reg_buffer[15], 15'b000000000010101)^gf_mul(reg_buffer[16], 15'b000000100000100)^gf_mul(reg_buffer[17], 15'b001010001010000)^gf_mul(reg_buffer[18], 15'b001010001000110);
	elp_eval[32]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000101000)^gf_mul(reg_buffer[2], 15'b000010001000000)^gf_mul(reg_buffer[3], 15'b010101000000011)^gf_mul(reg_buffer[4], 15'b001000001100000)^gf_mul(reg_buffer[5], 15'b000111100001111)^gf_mul(reg_buffer[6], 15'b001100110011101)^gf_mul(reg_buffer[7], 15'b111111101000001)^gf_mul(reg_buffer[8], 15'b001001000000000)^gf_mul(reg_buffer[9], 15'b101000000001111)^gf_mul(reg_buffer[10], 15'b000000110101011)^gf_mul(reg_buffer[11], 15'b011100000111000)^gf_mul(reg_buffer[12], 15'b100011011010111)^gf_mul(reg_buffer[13], 15'b110110001100111)^gf_mul(reg_buffer[14], 15'b110111111111111)^gf_mul(reg_buffer[15], 15'b000000000111111)^gf_mul(reg_buffer[16], 15'b000011000011000)^gf_mul(reg_buffer[17], 15'b111001111000011)^gf_mul(reg_buffer[18], 15'b110011001010101);
	elp_eval[33]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000001010000)^gf_mul(reg_buffer[2], 15'b001000100000000)^gf_mul(reg_buffer[3], 15'b101000000011110)^gf_mul(reg_buffer[4], 15'b000011000000110)^gf_mul(reg_buffer[5], 15'b110000111100101)^gf_mul(reg_buffer[6], 15'b110011101010100)^gf_mul(reg_buffer[7], 15'b010000000000001)^gf_mul(reg_buffer[8], 15'b000000001101100)^gf_mul(reg_buffer[9], 15'b001110111000000)^gf_mul(reg_buffer[10], 15'b010110000010111)^gf_mul(reg_buffer[11], 15'b100010010000101)^gf_mul(reg_buffer[12], 15'b110100101101110)^gf_mul(reg_buffer[13], 15'b100110100101011)^gf_mul(reg_buffer[14], 15'b001100000000001)^gf_mul(reg_buffer[15], 15'b000000001000001)^gf_mul(reg_buffer[16], 15'b001010001010000)^gf_mul(reg_buffer[17], 15'b101000100011000)^gf_mul(reg_buffer[18], 15'b101011111100110);
	elp_eval[34]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000010100000)^gf_mul(reg_buffer[2], 15'b100010000000000)^gf_mul(reg_buffer[3], 15'b000000011111111)^gf_mul(reg_buffer[4], 15'b110000001100000)^gf_mul(reg_buffer[5], 15'b011110010001000)^gf_mul(reg_buffer[6], 15'b101010101010101)^gf_mul(reg_buffer[7], 15'b000000011100000)^gf_mul(reg_buffer[8], 15'b110110000000000)^gf_mul(reg_buffer[9], 15'b000000010011001)^gf_mul(reg_buffer[10], 15'b101111110100000)^gf_mul(reg_buffer[11], 15'b010010011011000)^gf_mul(reg_buffer[12], 15'b111011101110111)^gf_mul(reg_buffer[13], 15'b101010111011110)^gf_mul(reg_buffer[14], 15'b101010000000000)^gf_mul(reg_buffer[15], 15'b000000011000011)^gf_mul(reg_buffer[16], 15'b111100111100000)^gf_mul(reg_buffer[17], 15'b100110010101001)^gf_mul(reg_buffer[18], 15'b100000101000001);
	elp_eval[35]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000101000000)^gf_mul(reg_buffer[2], 15'b001000000000110)^gf_mul(reg_buffer[3], 15'b000011111111000)^gf_mul(reg_buffer[4], 15'b000011000010100)^gf_mul(reg_buffer[5], 15'b001000100010001)^gf_mul(reg_buffer[6], 15'b101010100111110)^gf_mul(reg_buffer[7], 15'b111000000000000)^gf_mul(reg_buffer[8], 15'b000000101101000)^gf_mul(reg_buffer[9], 15'b011001000000110)^gf_mul(reg_buffer[10], 15'b000011100000111)^gf_mul(reg_buffer[11], 15'b100011011010111)^gf_mul(reg_buffer[12], 15'b110001100110010)^gf_mul(reg_buffer[13], 15'b111111110011001)^gf_mul(reg_buffer[14], 15'b111111000000000)^gf_mul(reg_buffer[15], 15'b000000101000101)^gf_mul(reg_buffer[16], 15'b001010001000110)^gf_mul(reg_buffer[17], 15'b101011111100110)^gf_mul(reg_buffer[18], 15'b001111000001100);
	elp_eval[36]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000001010000000)^gf_mul(reg_buffer[2], 15'b100000000011000)^gf_mul(reg_buffer[3], 15'b011111111000000)^gf_mul(reg_buffer[4], 15'b110000101000000)^gf_mul(reg_buffer[5], 15'b010001000101100)^gf_mul(reg_buffer[6], 15'b100111111111110)^gf_mul(reg_buffer[7], 15'b000000010010000)^gf_mul(reg_buffer[8], 15'b110100000000110)^gf_mul(reg_buffer[9], 15'b000110101011000)^gf_mul(reg_buffer[10], 15'b001110001001000)^gf_mul(reg_buffer[11], 15'b011010010110111)^gf_mul(reg_buffer[12], 15'b011010010101010)^gf_mul(reg_buffer[13], 15'b000000000101010)^gf_mul(reg_buffer[14], 15'b100000100000000)^gf_mul(reg_buffer[15], 15'b000001111001111)^gf_mul(reg_buffer[16], 15'b111100110010100)^gf_mul(reg_buffer[17], 15'b110000010100001)^gf_mul(reg_buffer[18], 15'b001000010100110);
	elp_eval[37]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000010100000000)^gf_mul(reg_buffer[2], 15'b000000001100110)^gf_mul(reg_buffer[3], 15'b111111000000101)^gf_mul(reg_buffer[4], 15'b001010000010100)^gf_mul(reg_buffer[5], 15'b100010110011000)^gf_mul(reg_buffer[6], 15'b111111111101001)^gf_mul(reg_buffer[7], 15'b100100000000000)^gf_mul(reg_buffer[8], 15'b000011101110000)^gf_mul(reg_buffer[9], 15'b011000001011111)^gf_mul(reg_buffer[10], 15'b010000100100110)^gf_mul(reg_buffer[11], 15'b011110111011101)^gf_mul(reg_buffer[12], 15'b010101110111111)^gf_mul(reg_buffer[13], 15'b100000000011110)^gf_mul(reg_buffer[14], 15'b110000110000000)^gf_mul(reg_buffer[15], 15'b000010001010001)^gf_mul(reg_buffer[16], 15'b001010101111110)^gf_mul(reg_buffer[17], 15'b000011110000011)^gf_mul(reg_buffer[18], 15'b000111101010101);
	elp_eval[38]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000101000000000)^gf_mul(reg_buffer[2], 15'b000000110011000)^gf_mul(reg_buffer[3], 15'b111000000100001)^gf_mul(reg_buffer[4], 15'b100000101000110)^gf_mul(reg_buffer[5], 15'b011001100110011)^gf_mul(reg_buffer[6], 15'b111101000000001)^gf_mul(reg_buffer[7], 15'b000000011011000)^gf_mul(reg_buffer[8], 15'b111000000010010)^gf_mul(reg_buffer[9], 15'b011111101000011)^gf_mul(reg_buffer[10], 15'b001101100011011)^gf_mul(reg_buffer[11], 15'b110110001100111)^gf_mul(reg_buffer[12], 15'b111111110011001)^gf_mul(reg_buffer[13], 15'b111000000001001)^gf_mul(reg_buffer[14], 15'b101000101000000)^gf_mul(reg_buffer[15], 15'b000110011110011)^gf_mul(reg_buffer[16], 15'b111111100000100)^gf_mul(reg_buffer[17], 15'b010001000010100)^gf_mul(reg_buffer[18], 15'b000111111111011);
	elp_eval[39]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b001010000000000)^gf_mul(reg_buffer[2], 15'b000011001100000)^gf_mul(reg_buffer[3], 15'b000000100000001)^gf_mul(reg_buffer[4], 15'b001010001111000)^gf_mul(reg_buffer[5], 15'b110011001110100)^gf_mul(reg_buffer[6], 15'b000000000000111)^gf_mul(reg_buffer[7], 15'b110110000000000)^gf_mul(reg_buffer[8], 15'b001001100100000)^gf_mul(reg_buffer[9], 15'b000011100000111)^gf_mul(reg_buffer[10], 15'b110110101101000)^gf_mul(reg_buffer[11], 15'b011001101001010)^gf_mul(reg_buffer[12], 15'b000000000010101)^gf_mul(reg_buffer[13], 15'b000010000000110)^gf_mul(reg_buffer[14], 15'b111100111100000)^gf_mul(reg_buffer[15], 15'b001010100010101)^gf_mul(reg_buffer[16], 15'b000001000011110)^gf_mul(reg_buffer[17], 15'b001100011110101)^gf_mul(reg_buffer[18], 15'b000000001101011);
	elp_eval[40]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b010100000000000)^gf_mul(reg_buffer[2], 15'b001100110000000)^gf_mul(reg_buffer[3], 15'b000100000001000)^gf_mul(reg_buffer[4], 15'b100011110000110)^gf_mul(reg_buffer[5], 15'b100111010101011)^gf_mul(reg_buffer[6], 15'b000000111000000)^gf_mul(reg_buffer[7], 15'b000000010110100)^gf_mul(reg_buffer[8], 15'b010000001101010)^gf_mul(reg_buffer[9], 15'b000111000100100)^gf_mul(reg_buffer[10], 15'b010010110111101)^gf_mul(reg_buffer[11], 15'b101010101011100)^gf_mul(reg_buffer[12], 15'b101000000000110)^gf_mul(reg_buffer[13], 15'b100001100000011)^gf_mul(reg_buffer[14], 15'b100010100010000)^gf_mul(reg_buffer[15], 15'b011111100111111)^gf_mul(reg_buffer[16], 15'b000110001000100)^gf_mul(reg_buffer[17], 15'b010010001111111)^gf_mul(reg_buffer[18], 15'b000010111101000);
	elp_eval[41]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b101000000000000)^gf_mul(reg_buffer[2], 15'b110011000000000)^gf_mul(reg_buffer[3], 15'b100000001000000)^gf_mul(reg_buffer[4], 15'b111100001111000)^gf_mul(reg_buffer[5], 15'b101010101010101)^gf_mul(reg_buffer[6], 15'b111000000000000)^gf_mul(reg_buffer[7], 15'b101101000000000)^gf_mul(reg_buffer[8], 15'b110101011000000)^gf_mul(reg_buffer[9], 15'b100100001001000)^gf_mul(reg_buffer[10], 15'b111011101110111)^gf_mul(reg_buffer[11], 15'b110111111111111)^gf_mul(reg_buffer[12], 15'b111111000000000)^gf_mul(reg_buffer[13], 15'b101000101000000)^gf_mul(reg_buffer[14], 15'b110011110011000)^gf_mul(reg_buffer[15], 15'b100000101000001)^gf_mul(reg_buffer[16], 15'b010100110011000)^gf_mul(reg_buffer[17], 15'b011001000000001)^gf_mul(reg_buffer[18], 15'b111000111000000);
	elp_eval[42]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b010000000000011)^gf_mul(reg_buffer[2], 15'b001100000000101)^gf_mul(reg_buffer[3], 15'b000001000001100)^gf_mul(reg_buffer[4], 15'b000011110010001)^gf_mul(reg_buffer[5], 15'b010101010011111)^gf_mul(reg_buffer[6], 15'b000000001001000)^gf_mul(reg_buffer[7], 15'b000000011101110)^gf_mul(reg_buffer[8], 15'b100000101111111)^gf_mul(reg_buffer[9], 15'b001001101100011)^gf_mul(reg_buffer[10], 15'b101100011001101)^gf_mul(reg_buffer[11], 15'b111001100000001)^gf_mul(reg_buffer[12], 15'b001000001000000)^gf_mul(reg_buffer[13], 15'b011110011110000)^gf_mul(reg_buffer[14], 15'b101010001010100)^gf_mul(reg_buffer[15], 15'b100001111000000)^gf_mul(reg_buffer[16], 15'b111010101010011)^gf_mul(reg_buffer[17], 15'b101100000001010)^gf_mul(reg_buffer[18], 15'b001001000011011);
	elp_eval[43]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b100000000000110)^gf_mul(reg_buffer[2], 15'b110000000010100)^gf_mul(reg_buffer[3], 15'b001000001100000)^gf_mul(reg_buffer[4], 15'b111100100010000)^gf_mul(reg_buffer[5], 15'b101001111111110)^gf_mul(reg_buffer[6], 15'b001001000000000)^gf_mul(reg_buffer[7], 15'b111011100000000)^gf_mul(reg_buffer[8], 15'b111111010000110)^gf_mul(reg_buffer[9], 15'b100011011010111)^gf_mul(reg_buffer[10], 15'b011001101001010)^gf_mul(reg_buffer[11], 15'b000000101010000)^gf_mul(reg_buffer[12], 15'b000011000011000)^gf_mul(reg_buffer[13], 15'b001000101000100)^gf_mul(reg_buffer[14], 15'b111111001111110)^gf_mul(reg_buffer[15], 15'b100010001000011)^gf_mul(reg_buffer[16], 15'b011111111101100)^gf_mul(reg_buffer[17], 15'b010000001110001)^gf_mul(reg_buffer[18], 15'b011000101101101);
	elp_eval[44]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000001111)^gf_mul(reg_buffer[2], 15'b000000001010101)^gf_mul(reg_buffer[3], 15'b000001100000011)^gf_mul(reg_buffer[4], 15'b001000100010001)^gf_mul(reg_buffer[5], 15'b111111111111100)^gf_mul(reg_buffer[6], 15'b000000000011011)^gf_mul(reg_buffer[7], 15'b000000010011001)^gf_mul(reg_buffer[8], 15'b000011100000111)^gf_mul(reg_buffer[9], 15'b010110100101101)^gf_mul(reg_buffer[10], 15'b010101010101110)^gf_mul(reg_buffer[11], 15'b000000000111111)^gf_mul(reg_buffer[12], 15'b000000101000101)^gf_mul(reg_buffer[13], 15'b000110011110011)^gf_mul(reg_buffer[14], 15'b100000101000001)^gf_mul(reg_buffer[15], 15'b100110011000110)^gf_mul(reg_buffer[16], 15'b000000001101011)^gf_mul(reg_buffer[17], 15'b000001001001001)^gf_mul(reg_buffer[18], 15'b001110110110111);
	elp_eval[45]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000011110)^gf_mul(reg_buffer[2], 15'b000000101010100)^gf_mul(reg_buffer[3], 15'b001100000011000)^gf_mul(reg_buffer[4], 15'b001000100010110)^gf_mul(reg_buffer[5], 15'b111111110100001)^gf_mul(reg_buffer[6], 15'b000011011000000)^gf_mul(reg_buffer[7], 15'b100110010000000)^gf_mul(reg_buffer[8], 15'b000011100010010)^gf_mul(reg_buffer[9], 15'b101101111011100)^gf_mul(reg_buffer[10], 15'b011101111111111)^gf_mul(reg_buffer[11], 15'b111100000000101)^gf_mul(reg_buffer[12], 15'b101000001111000)^gf_mul(reg_buffer[13], 15'b110010101000100)^gf_mul(reg_buffer[14], 15'b010000111100000)^gf_mul(reg_buffer[15], 15'b101010101001001)^gf_mul(reg_buffer[16], 15'b000000101111010)^gf_mul(reg_buffer[17], 15'b001101101101100)^gf_mul(reg_buffer[18], 15'b011011011001110);
	elp_eval[46]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000111100)^gf_mul(reg_buffer[2], 15'b000010101010000)^gf_mul(reg_buffer[3], 15'b100000011000011)^gf_mul(reg_buffer[4], 15'b001000101100110)^gf_mul(reg_buffer[5], 15'b111010000000001)^gf_mul(reg_buffer[6], 15'b011000000000101)^gf_mul(reg_buffer[7], 15'b100000011010100)^gf_mul(reg_buffer[8], 15'b001001000010010)^gf_mul(reg_buffer[9], 15'b011101110110001)^gf_mul(reg_buffer[10], 15'b111111001100001)^gf_mul(reg_buffer[11], 15'b010000010000000)^gf_mul(reg_buffer[12], 15'b001111000010001)^gf_mul(reg_buffer[13], 15'b010101111110011)^gf_mul(reg_buffer[14], 15'b011000100010000)^gf_mul(reg_buffer[15], 15'b111111111011000)^gf_mul(reg_buffer[16], 15'b000011100011100)^gf_mul(reg_buffer[17], 15'b011011011010011)^gf_mul(reg_buffer[18], 15'b101101010011111);
	elp_eval[47]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000001111000)^gf_mul(reg_buffer[2], 15'b001010101000000)^gf_mul(reg_buffer[3], 15'b000011000010100)^gf_mul(reg_buffer[4], 15'b001011001100110)^gf_mul(reg_buffer[5], 15'b000000000000111)^gf_mul(reg_buffer[6], 15'b000000101101000)^gf_mul(reg_buffer[7], 15'b110101011000000)^gf_mul(reg_buffer[8], 15'b001001001101100)^gf_mul(reg_buffer[9], 15'b110001100110010)^gf_mul(reg_buffer[10], 15'b000000000010101)^gf_mul(reg_buffer[11], 15'b000011000011000)^gf_mul(reg_buffer[12], 15'b001010001000110)^gf_mul(reg_buffer[13], 15'b111111100000100)^gf_mul(reg_buffer[14], 15'b010100110011000)^gf_mul(reg_buffer[15], 15'b000000001101011)^gf_mul(reg_buffer[16], 15'b001001001001000)^gf_mul(reg_buffer[17], 15'b110110111010010)^gf_mul(reg_buffer[18], 15'b111110100011010);
	elp_eval[48]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000011110000)^gf_mul(reg_buffer[2], 15'b101010100000000)^gf_mul(reg_buffer[3], 15'b011000010100000)^gf_mul(reg_buffer[4], 15'b110011001100110)^gf_mul(reg_buffer[5], 15'b000000011100000)^gf_mul(reg_buffer[6], 15'b101101000000000)^gf_mul(reg_buffer[7], 15'b110000010111110)^gf_mul(reg_buffer[8], 15'b110110001101100)^gf_mul(reg_buffer[9], 15'b110011010010100)^gf_mul(reg_buffer[10], 15'b101010000000000)^gf_mul(reg_buffer[11], 15'b100000010100011)^gf_mul(reg_buffer[12], 15'b110011110011000)^gf_mul(reg_buffer[13], 15'b010000001000011)^gf_mul(reg_buffer[14], 15'b011110101010100)^gf_mul(reg_buffer[15], 15'b000000010111101)^gf_mul(reg_buffer[16], 15'b110110110110000)^gf_mul(reg_buffer[17], 15'b101100111010111)^gf_mul(reg_buffer[18], 15'b011100101101000);
	elp_eval[49]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000111100000)^gf_mul(reg_buffer[2], 15'b101010000000110)^gf_mul(reg_buffer[3], 15'b000010100000101)^gf_mul(reg_buffer[4], 15'b110011001110100)^gf_mul(reg_buffer[5], 15'b001110000000000)^gf_mul(reg_buffer[6], 15'b000000001110111)^gf_mul(reg_buffer[7], 15'b101111110100000)^gf_mul(reg_buffer[8], 15'b110110101101000)^gf_mul(reg_buffer[9], 15'b010101010101110)^gf_mul(reg_buffer[10], 15'b000011111100000)^gf_mul(reg_buffer[11], 15'b001010000011110)^gf_mul(reg_buffer[12], 15'b001010100010101)^gf_mul(reg_buffer[13], 15'b111100000110000)^gf_mul(reg_buffer[14], 15'b010001111111110)^gf_mul(reg_buffer[15], 15'b000000111000111)^gf_mul(reg_buffer[16], 15'b110110110100110)^gf_mul(reg_buffer[17], 15'b010100111101101)^gf_mul(reg_buffer[18], 15'b101110111001100);
	elp_eval[50]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000001111000000)^gf_mul(reg_buffer[2], 15'b101000000011110)^gf_mul(reg_buffer[3], 15'b010100000101000)^gf_mul(reg_buffer[4], 15'b110011101010100)^gf_mul(reg_buffer[5], 15'b000000000001001)^gf_mul(reg_buffer[6], 15'b001110111000000)^gf_mul(reg_buffer[7], 15'b101000011100001)^gf_mul(reg_buffer[8], 15'b110100101101110)^gf_mul(reg_buffer[9], 15'b101110111111110)^gf_mul(reg_buffer[10], 15'b000000001000001)^gf_mul(reg_buffer[11], 15'b111001111000011)^gf_mul(reg_buffer[12], 15'b101011111100110)^gf_mul(reg_buffer[13], 15'b010001000010100)^gf_mul(reg_buffer[14], 15'b011001000000001)^gf_mul(reg_buffer[15], 15'b000001001001001)^gf_mul(reg_buffer[16], 15'b110110111010010)^gf_mul(reg_buffer[17], 15'b110100011011001)^gf_mul(reg_buffer[18], 15'b011001010110010);
	elp_eval[51]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000011110000000)^gf_mul(reg_buffer[2], 15'b100000001111110)^gf_mul(reg_buffer[3], 15'b100000101000110)^gf_mul(reg_buffer[4], 15'b111010101010100)^gf_mul(reg_buffer[5], 15'b000000100100000)^gf_mul(reg_buffer[6], 15'b111000000010010)^gf_mul(reg_buffer[7], 15'b111000001110000)^gf_mul(reg_buffer[8], 15'b110111101110110)^gf_mul(reg_buffer[9], 15'b111111110011001)^gf_mul(reg_buffer[10], 15'b000010000000110)^gf_mul(reg_buffer[11], 15'b001000101000100)^gf_mul(reg_buffer[12], 15'b111111100000100)^gf_mul(reg_buffer[13], 15'b001100110001111)^gf_mul(reg_buffer[14], 15'b110101100000000)^gf_mul(reg_buffer[15], 15'b000011011011011)^gf_mul(reg_buffer[16], 15'b110110011101010)^gf_mul(reg_buffer[17], 15'b110010110100011)^gf_mul(reg_buffer[18], 15'b011111010111111);
	elp_eval[52]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000111100000000)^gf_mul(reg_buffer[2], 15'b000000111111110)^gf_mul(reg_buffer[3], 15'b000101000111100)^gf_mul(reg_buffer[4], 15'b101010101010010)^gf_mul(reg_buffer[5], 15'b010010000000000)^gf_mul(reg_buffer[6], 15'b000010011001000)^gf_mul(reg_buffer[7], 15'b011100010010000)^gf_mul(reg_buffer[8], 15'b111011101100010)^gf_mul(reg_buffer[9], 15'b011000000000010)^gf_mul(reg_buffer[10], 15'b001100001100000)^gf_mul(reg_buffer[11], 15'b010001100111100)^gf_mul(reg_buffer[12], 15'b101000000100000)^gf_mul(reg_buffer[13], 15'b110101010100101)^gf_mul(reg_buffer[14], 15'b101111010000000)^gf_mul(reg_buffer[15], 15'b000101101101101)^gf_mul(reg_buffer[16], 15'b110101001111010)^gf_mul(reg_buffer[17], 15'b011101110011011)^gf_mul(reg_buffer[18], 15'b001111000000100);
	elp_eval[53]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b001111000000000)^gf_mul(reg_buffer[2], 15'b000011111111000)^gf_mul(reg_buffer[3], 15'b101000111100000)^gf_mul(reg_buffer[4], 15'b101010100111110)^gf_mul(reg_buffer[5], 15'b000000000011011)^gf_mul(reg_buffer[6], 15'b011001000000110)^gf_mul(reg_buffer[7], 15'b100100001001000)^gf_mul(reg_buffer[8], 15'b110001100110010)^gf_mul(reg_buffer[9], 15'b000010101000000)^gf_mul(reg_buffer[10], 15'b000000101000101)^gf_mul(reg_buffer[11], 15'b110011001010101)^gf_mul(reg_buffer[12], 15'b001111000001100)^gf_mul(reg_buffer[13], 15'b000111111111011)^gf_mul(reg_buffer[14], 15'b111000111000000)^gf_mul(reg_buffer[15], 15'b001110110110111)^gf_mul(reg_buffer[16], 15'b111110100011010)^gf_mul(reg_buffer[17], 15'b011001010110010)^gf_mul(reg_buffer[18], 15'b001000001100110);
	elp_eval[54]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b011110000000000)^gf_mul(reg_buffer[2], 15'b001111111100000)^gf_mul(reg_buffer[3], 15'b000111100001111)^gf_mul(reg_buffer[4], 15'b101001111111110)^gf_mul(reg_buffer[5], 15'b000001101100000)^gf_mul(reg_buffer[6], 15'b000000110101011)^gf_mul(reg_buffer[7], 15'b010010011011000)^gf_mul(reg_buffer[8], 15'b011001101001010)^gf_mul(reg_buffer[9], 15'b000000000111111)^gf_mul(reg_buffer[10], 15'b001010000011110)^gf_mul(reg_buffer[11], 15'b010001010101111)^gf_mul(reg_buffer[12], 15'b100010001000011)^gf_mul(reg_buffer[13], 15'b110010000000010)^gf_mul(reg_buffer[14], 15'b100100100100000)^gf_mul(reg_buffer[15], 15'b010011011011001)^gf_mul(reg_buffer[16], 15'b000111001011010)^gf_mul(reg_buffer[17], 15'b101111101011110)^gf_mul(reg_buffer[18], 15'b000010101010101);
	elp_eval[55]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b111100000000000)^gf_mul(reg_buffer[2], 15'b111111110000000)^gf_mul(reg_buffer[3], 15'b111100001111000)^gf_mul(reg_buffer[4], 15'b011111111111110)^gf_mul(reg_buffer[5], 15'b110110000000000)^gf_mul(reg_buffer[6], 15'b110101011000000)^gf_mul(reg_buffer[7], 15'b110110001101100)^gf_mul(reg_buffer[8], 15'b100101010101010)^gf_mul(reg_buffer[9], 15'b111111000000000)^gf_mul(reg_buffer[10], 15'b111100111100000)^gf_mul(reg_buffer[11], 15'b111111001111110)^gf_mul(reg_buffer[12], 15'b010100110011000)^gf_mul(reg_buffer[13], 15'b110101100000000)^gf_mul(reg_buffer[14], 15'b110110110110000)^gf_mul(reg_buffer[15], 15'b110101101101011)^gf_mul(reg_buffer[16], 15'b010010111011100)^gf_mul(reg_buffer[17], 15'b000011110000001)^gf_mul(reg_buffer[18], 15'b111111111111000);
	elp_eval[56]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b111000000000011)^gf_mul(reg_buffer[2], 15'b111111000000101)^gf_mul(reg_buffer[3], 15'b100001111001001)^gf_mul(reg_buffer[4], 15'b111111111101001)^gf_mul(reg_buffer[5], 15'b000000000101101)^gf_mul(reg_buffer[6], 15'b011000001011111)^gf_mul(reg_buffer[7], 15'b011011010110100)^gf_mul(reg_buffer[8], 15'b010101110111111)^gf_mul(reg_buffer[9], 15'b000001000001000)^gf_mul(reg_buffer[10], 15'b000010001010001)^gf_mul(reg_buffer[11], 15'b111100000101001)^gf_mul(reg_buffer[12], 15'b000111101010101)^gf_mul(reg_buffer[13], 15'b010111101000000)^gf_mul(reg_buffer[14], 15'b101101101101000)^gf_mul(reg_buffer[15], 15'b011110110111110)^gf_mul(reg_buffer[16], 15'b101110011001011)^gf_mul(reg_buffer[17], 15'b010001000001100)^gf_mul(reg_buffer[18], 15'b000000001011000);
	elp_eval[57]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b110000000000101)^gf_mul(reg_buffer[2], 15'b111100000010001)^gf_mul(reg_buffer[3], 15'b001111001000100)^gf_mul(reg_buffer[4], 15'b111111010000001)^gf_mul(reg_buffer[5], 15'b000010110100000)^gf_mul(reg_buffer[6], 15'b001011111101000)^gf_mul(reg_buffer[7], 15'b101101001011010)^gf_mul(reg_buffer[8], 15'b011111111111001)^gf_mul(reg_buffer[9], 15'b001000000011000)^gf_mul(reg_buffer[10], 15'b100010001100110)^gf_mul(reg_buffer[11], 15'b100000010000110)^gf_mul(reg_buffer[12], 15'b101001000111110)^gf_mul(reg_buffer[13], 15'b001110001110000)^gf_mul(reg_buffer[14], 15'b111011011011100)^gf_mul(reg_buffer[15], 15'b100011011000010)^gf_mul(reg_buffer[16], 15'b100101010111111)^gf_mul(reg_buffer[17], 15'b001100001010101)^gf_mul(reg_buffer[18], 15'b000011101000000);
	elp_eval[58]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b100000000001001)^gf_mul(reg_buffer[2], 15'b110000001000001)^gf_mul(reg_buffer[3], 15'b111001000100011)^gf_mul(reg_buffer[4], 15'b110100000000001)^gf_mul(reg_buffer[5], 15'b011010000000011)^gf_mul(reg_buffer[6], 15'b111101000011101)^gf_mul(reg_buffer[7], 15'b010110111101110)^gf_mul(reg_buffer[8], 15'b111100110000001)^gf_mul(reg_buffer[9], 15'b011000011000000)^gf_mul(reg_buffer[10], 15'b001111001100101)^gf_mul(reg_buffer[11], 15'b011110000011000)^gf_mul(reg_buffer[12], 15'b111111011001001)^gf_mul(reg_buffer[13], 15'b000100100100100)^gf_mul(reg_buffer[14], 15'b100110110110010)^gf_mul(reg_buffer[15], 15'b100101101000101)^gf_mul(reg_buffer[16], 15'b011111110000111)^gf_mul(reg_buffer[17], 15'b010001111111111)^gf_mul(reg_buffer[18], 15'b100111000000000);
	elp_eval[59]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000010001)^gf_mul(reg_buffer[2], 15'b000000100000001)^gf_mul(reg_buffer[3], 15'b001000100010001)^gf_mul(reg_buffer[4], 15'b000000000000111)^gf_mul(reg_buffer[5], 15'b000000001110111)^gf_mul(reg_buffer[6], 15'b000011100000111)^gf_mul(reg_buffer[7], 15'b111011101110111)^gf_mul(reg_buffer[8], 15'b000000000010101)^gf_mul(reg_buffer[9], 15'b000000101000101)^gf_mul(reg_buffer[10], 15'b001010100010101)^gf_mul(reg_buffer[11], 15'b100010001000011)^gf_mul(reg_buffer[12], 15'b000000001101011)^gf_mul(reg_buffer[13], 15'b000011011011011)^gf_mul(reg_buffer[14], 15'b110101101101011)^gf_mul(reg_buffer[15], 15'b101110111001100)^gf_mul(reg_buffer[16], 15'b000000100010001)^gf_mul(reg_buffer[17], 15'b001000000000001)^gf_mul(reg_buffer[18], 15'b001000000010111);
	elp_eval[60]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000000100010)^gf_mul(reg_buffer[2], 15'b000010000000100)^gf_mul(reg_buffer[3], 15'b000100010001011)^gf_mul(reg_buffer[4], 15'b000000001110000)^gf_mul(reg_buffer[5], 15'b000111011100000)^gf_mul(reg_buffer[6], 15'b100000111000101)^gf_mul(reg_buffer[7], 15'b011101100011001)^gf_mul(reg_buffer[8], 15'b001010100000000)^gf_mul(reg_buffer[9], 15'b000101000001111)^gf_mul(reg_buffer[10], 15'b101010111111000)^gf_mul(reg_buffer[11], 15'b001010011001100)^gf_mul(reg_buffer[12], 15'b011000000010111)^gf_mul(reg_buffer[13], 15'b110001011011010)^gf_mul(reg_buffer[14], 15'b001111011011111)^gf_mul(reg_buffer[15], 15'b110011001010111)^gf_mul(reg_buffer[16], 15'b000011001100110)^gf_mul(reg_buffer[17], 15'b100000000001111)^gf_mul(reg_buffer[18], 15'b000000111001101);
	elp_eval[61]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000001000100)^gf_mul(reg_buffer[2], 15'b001000000010000)^gf_mul(reg_buffer[3], 15'b100010001011000)^gf_mul(reg_buffer[4], 15'b000011100000000)^gf_mul(reg_buffer[5], 15'b101110000000101)^gf_mul(reg_buffer[6], 15'b111000100100000)^gf_mul(reg_buffer[7], 15'b000110011001101)^gf_mul(reg_buffer[8], 15'b000000001111110)^gf_mul(reg_buffer[9], 15'b001111001111000)^gf_mul(reg_buffer[10], 15'b110011111110001)^gf_mul(reg_buffer[11], 15'b110001111010100)^gf_mul(reg_buffer[12], 15'b111101000000110)^gf_mul(reg_buffer[13], 15'b110100111011010)^gf_mul(reg_buffer[14], 15'b101000110110001)^gf_mul(reg_buffer[15], 15'b010101011111010)^gf_mul(reg_buffer[16], 15'b001010101010100)^gf_mul(reg_buffer[17], 15'b000000001001110)^gf_mul(reg_buffer[18], 15'b001001010111000);
	elp_eval[62]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000010001000)^gf_mul(reg_buffer[2], 15'b100000001000000)^gf_mul(reg_buffer[3], 15'b010001011001100)^gf_mul(reg_buffer[4], 15'b111000000000000)^gf_mul(reg_buffer[5], 15'b000000010011001)^gf_mul(reg_buffer[6], 15'b100100001001000)^gf_mul(reg_buffer[7], 15'b110011010010100)^gf_mul(reg_buffer[8], 15'b111111000000000)^gf_mul(reg_buffer[9], 15'b111000010001011)^gf_mul(reg_buffer[10], 15'b100000101000001)^gf_mul(reg_buffer[11], 15'b010101001000111)^gf_mul(reg_buffer[12], 15'b111000111000000)^gf_mul(reg_buffer[13], 15'b110111010011010)^gf_mul(reg_buffer[14], 15'b011100101101000)^gf_mul(reg_buffer[15], 15'b111111100001110)^gf_mul(reg_buffer[16], 15'b111111111111000)^gf_mul(reg_buffer[17], 15'b000001101001000)^gf_mul(reg_buffer[18], 15'b011111001000101);
	elp_eval[63]=	reg_buffer[0]^gf_mul(reg_buffer[1], 15'b000000100010000)^gf_mul(reg_buffer[2], 15'b000000100000110)^gf_mul(reg_buffer[3], 15'b001011001100110)^gf_mul(reg_buffer[4], 15'b000000000010010)^gf_mul(reg_buffer[5], 15'b001001100100000)^gf_mul(reg_buffer[6], 15'b001001001101100)^gf_mul(reg_buffer[7], 15'b100101010101010)^gf_mul(reg_buffer[8], 15'b000000100000100)^gf_mul(reg_buffer[9], 15'b001010001000110)^gf_mul(reg_buffer[10], 15'b000001000011110)^gf_mul(reg_buffer[11], 15'b011111111101100)^gf_mul(reg_buffer[12], 15'b001001001001000)^gf_mul(reg_buffer[13], 15'b110110011101010)^gf_mul(reg_buffer[14], 15'b010010111011100)^gf_mul(reg_buffer[15], 15'b000000100010001)^gf_mul(reg_buffer[16], 15'b000000000010110)^gf_mul(reg_buffer[17], 15'b001011101100000)^gf_mul(reg_buffer[18], 15'b001011001110100);
	return elp_eval;
endfunction

(* noinline *)
function Vector#(19, Bit#(15)) update_reg_buffer(Vector#(19, Bit#(15)) reg_buffer);
	Vector#(19, Bit#(15)) reg_buffer_updated;
	reg_buffer_updated[0] = 	reg_buffer[0];
	reg_buffer_updated[1] = 	gf_mul(reg_buffer[1], 15'b000000100010000);
	reg_buffer_updated[2] = 	gf_mul(reg_buffer[2], 15'b000000100000110);
	reg_buffer_updated[3] = 	gf_mul(reg_buffer[3], 15'b001011001100110);
	reg_buffer_updated[4] = 	gf_mul(reg_buffer[4], 15'b000000000010010);
	reg_buffer_updated[5] = 	gf_mul(reg_buffer[5], 15'b001001100100000);
	reg_buffer_updated[6] = 	gf_mul(reg_buffer[6], 15'b001001001101100);
	reg_buffer_updated[7] = 	gf_mul(reg_buffer[7], 15'b100101010101010);
	reg_buffer_updated[8] = 	gf_mul(reg_buffer[8], 15'b000000100000100);
	reg_buffer_updated[9] = 	gf_mul(reg_buffer[9], 15'b001010001000110);
	reg_buffer_updated[10] = 	gf_mul(reg_buffer[10], 15'b000001000011110);
	reg_buffer_updated[11] = 	gf_mul(reg_buffer[11], 15'b011111111101100);
	reg_buffer_updated[12] = 	gf_mul(reg_buffer[12], 15'b001001001001000);
	reg_buffer_updated[13] = 	gf_mul(reg_buffer[13], 15'b110110011101010);
	reg_buffer_updated[14] = 	gf_mul(reg_buffer[14], 15'b010010111011100);
	reg_buffer_updated[15] = 	gf_mul(reg_buffer[15], 15'b000000100010001);
	reg_buffer_updated[16] = 	gf_mul(reg_buffer[16], 15'b000000000010110);
	reg_buffer_updated[17] = 	gf_mul(reg_buffer[17], 15'b001011101100000);
	reg_buffer_updated[18] = 	gf_mul(reg_buffer[18], 15'b001011001110100);
	return reg_buffer_updated;
endfunction

(* noinline *)
function Vector#(19, Bit#(15)) init_reg_buffer(Vector#(19, Bit#(15)) reg_buffer);
	Vector#(19, Bit#(15)) reg_init;
	reg_init[0] = 	reg_buffer[0];
	reg_init[1] = 	gf_mul(reg_buffer[1], 15'b010000010100111);
	reg_init[2] = 	gf_mul(reg_buffer[2], 15'b101110000010101);
	reg_init[3] = 	gf_mul(reg_buffer[3], 15'b000010110011100);
	reg_init[4] = 	gf_mul(reg_buffer[4], 15'b110011011110001);
	reg_init[5] = 	gf_mul(reg_buffer[5], 15'b001110000110100);
	reg_init[6] = 	gf_mul(reg_buffer[6], 15'b100000100110110);
	reg_init[7] = 	gf_mul(reg_buffer[7], 15'b000101001100011);
	reg_init[8] = 	gf_mul(reg_buffer[8], 15'b010110101111001);
	reg_init[9] = 	gf_mul(reg_buffer[9], 15'b110110001000100);
	reg_init[10] = 	gf_mul(reg_buffer[10], 15'b000001011110000);
	reg_init[11] = 	gf_mul(reg_buffer[11], 15'b010101100010010);
	reg_init[12] = 	gf_mul(reg_buffer[12], 15'b110010100010010);
	reg_init[13] = 	gf_mul(reg_buffer[13], 15'b111101101110000);
	reg_init[14] = 	gf_mul(reg_buffer[14], 15'b001010110011101);
	reg_init[15] = 	gf_mul(reg_buffer[15], 15'b011101001101010);
	reg_init[16] = 	gf_mul(reg_buffer[16], 15'b000110010100111);
	reg_init[17] = 	gf_mul(reg_buffer[17], 15'b000010101111111);
	reg_init[18] = 	gf_mul(reg_buffer[18], 15'b110100111110000);
	return reg_init;
endfunction


`include "encoder_logic_N16654_K16384.bsv"
`include "syndrome_logic_N16654_K16384.bsv"

endpackage: BCH_common

