function Bit#(32) get_output(UInt#(10) counter, UInt#(3) page_num);
	Bit#(32) enc_output = case (page_num)
		3'd0: get_output_page0(counter);
		3'd1: get_output_page1(counter);
		3'd2: get_output_page2(counter);
		3'd3: get_output_page3(counter);
		3'd4: get_output_page4(counter);
		3'd5: get_output_page5(counter);
		3'd6: get_output_page6(counter);
	endcase;
	return enc_output;
endfunction

function Bit#(32) get_output_page0(UInt#(10) counter);
	Bit#(32) out = case(counter)
		10'd0: 32'b00000000100000000000000000000000;
		10'd1: 32'b00000000000100000000000000000000;
		10'd2: 32'b00000000000000000000000000100000;
		10'd3: 32'b00000001000000000000000000010000;
		10'd4: 32'b00000100000000000000000000000000;
		10'd5: 32'b10000000000000000000000000000000;
		10'd6: 32'b00000000000000000000000100010000;
		10'd7: 32'b00000000000000000000000100000010;
		10'd8: 32'b00000000000000000000000100000010;
		10'd9: 32'b00000000000000000000000000000101;
		10'd10: 32'b00000001000000000000000000000100;
		10'd11: 32'b00000001000000000000000000010000;
		10'd12: 32'b00000000000100000000000000000000;
		10'd13: 32'b00000000001000000000000000000000;
		10'd14: 32'b00000000000000000000010000000000;
		10'd15: 32'b01000000000000000000000000000000;
		10'd16: 32'b00010000000000000000000000000010;
		10'd17: 32'b00000000000000000100000000000010;
		10'd18: 32'b00000000000000010000000000000001;
		10'd19: 32'b00000000000000000001000000000100;
		10'd20: 32'b00000000000000000000000000000011;
		10'd21: 32'b00000000000000010000000000000100;
		10'd22: 32'b00000000000000010000000000010000;
		10'd23: 32'b00100000000000000000000000000000;
		10'd24: 32'b00000000000000000100000000000000;
		10'd25: 32'b00000000000000000000000000000000;
		10'd26: 32'b00000000000000000000000000010000;
		10'd27: 32'b00000000000000000000000100000010;
		10'd28: 32'b00000001000000000000000000000100;
		10'd29: 32'b00000000000000000001000000000000;
		10'd30: 32'b00000000000000000000000000000010;
		10'd31: 32'b00000000000000001000000000000000;
		10'd32: 32'b00000000000000001000000000000000;
		10'd33: 32'b00000000010000000000000000000000;
		10'd34: 32'b00000000000000000100000000000010;
		10'd35: 32'b00000001000000000000000000000100;
		10'd36: 32'b01000000000000000000000000000010;
		10'd37: 32'b00000000010000000000000000000000;
		10'd38: 32'b00000000000000000001000000000100;
		10'd39: 32'b00100000000000000000000000000000;
		10'd40: 32'b00000000000000010000000000000010;
		10'd41: 32'b00000000000000010000000000000010;
		10'd42: 32'b00000000000100000000000000000100;
		10'd43: 32'b00000000000000000010000000000000;
		10'd44: 32'b00000000000000000000000100000001;
		10'd45: 32'b00000000000000000000001000000000;
		10'd46: 32'b00000000010000000000000000000000;
		10'd47: 32'b00000000000000000000000000100000;
		10'd48: 32'b00000000000000000000000000010000;
		10'd49: 32'b00000000000001000000000000000000;
		10'd50: 32'b00010000000000000000000000000010;
		10'd51: 32'b00000000000000000100000000000000;
		10'd52: 32'b00000000000000001000000000000000;
		10'd53: 32'b00000000000000000000000000000010;
		10'd54: 32'b01000000000000000000000000000010;
		10'd55: 32'b00001000000000000000000000000000;
		10'd56: 32'b00000000000000000000000000010100;
		10'd57: 32'b00000000000000000000000100000001;
		10'd58: 32'b00000000000000000000000001000000;
		10'd59: 32'b00000000000000000000000000000110;
		10'd60: 32'b00000000000000000000000100000010;
		10'd61: 32'b00000000000000000000000010000000;
		10'd62: 32'b00000000000000010000000000000000;
		10'd63: 32'b01000011000000011010000100001000;
		10'd64: 32'b00001000010000000000010000000000;
		10'd65: 32'b00000000000010001000000000000000;
		10'd66: 32'b01101001000001000000000001000000;
		10'd67: 32'b10000000000100010000000001000000;
		10'd68: 32'b00000000000000000000000010000000;
		10'd69: 32'b00000000100000000000000000000000;
		10'd70: 32'b00000100000000011001000000101010;
		10'd71: 32'b00100000000000000001000000000001;
		10'd72: 32'b00000100000110000000110000100010;
		10'd73: 32'b00000000000000000000000100000000;
		10'd74: 32'b01000000000000000000000000000000;
		10'd75: 32'b00000100000000000000000110000000;
		10'd76: 32'b00000000000000010000000000000000;
		10'd77: 32'b10000000000000000000001101010000;
		10'd78: 32'b00100000001001100000001000100100;
		10'd79: 32'b00000000010000001010011001010000;
		10'd80: 32'b00000000000000001000010000000000;
		10'd81: 32'b00000100010000000000100001000000;
		10'd82: 32'b00000001010000000010001000000000;
		10'd83: 32'b00000000000000000000000000110000;
		10'd84: 32'b00000000000000000001000100000000;
		10'd85: 32'b10000000000000000000010000000000;
		10'd86: 32'b00000000000000000000000000000010;
		10'd87: 32'b00000000000001010000000010000001;
		10'd88: 32'b00000100100001000100000101010000;
		10'd89: 32'b00000010000011000010001010000000;
		10'd90: 32'b00010000000001000010001000000000;
		10'd91: 32'b00000000000010000000010000000000;
		10'd92: 32'b00000100010000000000000001000000;
		10'd93: 32'b00000000000100000000010000000000;
		10'd94: 32'b00000010000000000000010100000010;
		10'd95: 32'b01000100000100000000000011000000;
		10'd96: 32'b00000000000000010000000000000000;
		10'd97: 32'b10001010000000001000000010000000;
		10'd98: 32'b00010000000000000000001000000000;
		10'd99: 32'b00000000000000000010010000000000;
		10'd100: 32'b01000000000000000100000000000000;
		10'd101: 32'b01000000000000000000000000001000;
		10'd102: 32'b00100000000000010000000001000001;
		10'd103: 32'b00000000000000000010000000000000;
		10'd104: 32'b00000010010100000110000100000000;
		10'd105: 32'b00000010010101001000000000010000;
		10'd106: 32'b00000000000000000100100000000011;
		10'd107: 32'b00101000100000100000000100000000;
		10'd108: 32'b00000010000000010000000000001000;
		10'd109: 32'b00000000001000100000000100000001;
		10'd110: 32'b00000000000000000000001000100000;
		10'd111: 32'b00000000000001100000010000000000;
		10'd112: 32'b10100000000001000100000000000001;
		10'd113: 32'b00000000000000000111100000010000;
		10'd114: 32'b10100000000001000000100000100000;
		10'd115: 32'b00100100000000001000000000000000;
		10'd116: 32'b01000010000000001000010000000000;
		10'd117: 32'b00001000000000000000001000000100;
		10'd118: 32'b00000000000000000000100000000010;
		10'd119: 32'b00000000010000100001000001000000;
		10'd120: 32'b00010100000000000001000000000010;
		10'd121: 32'b01100100000000000000000000011011;
		10'd122: 32'b00000000010000000001000000000001;
		10'd123: 32'b00100000000000000000001010000010;
		10'd124: 32'b00000000010000010000000000000100;
		10'd125: 32'b00000000001010000000000000000000;
		10'd126: 32'b00001001000000010100100000100010;
		10'd127: 32'b00000000000000000100000100000001;
		10'd128: 32'b00100000000000011000000000000010;
		10'd129: 32'b00000000000001000011000000011100;
		10'd130: 32'b00000000000000100000000010000010;
		10'd131: 32'b00000100000000000000000001110000;
		10'd132: 32'b00001000000000000000100010000010;
		10'd133: 32'b00000000101010000000000000000000;
		10'd134: 32'b01001010010000000001100000010000;
		10'd135: 32'b00101000001000000000000010100000;
		10'd136: 32'b00000000000000000000000000000000;
		10'd137: 32'b00000100000000001000000000000101;
		10'd138: 32'b10010000100001000000100000000000;
		10'd139: 32'b00000000000000000000110000000000;
		10'd140: 32'b00001000000000000000001100000000;
		10'd141: 32'b00010010000000000000011000001100;
		10'd142: 32'b00000010000001000001001000000000;
		10'd143: 32'b00000100000000010100000000000000;
		10'd144: 32'b01000000000001000000000000001000;
		10'd145: 32'b00000000000000000000000000000000;
		10'd146: 32'b01100100000010101000000000000000;
		10'd147: 32'b00100100001010000100000000000001;
		10'd148: 32'b00000000000100000100000000000000;
		10'd149: 32'b00100000000000000100000001000000;
		10'd150: 32'b00000000100000000000100011000000;
		10'd151: 32'b00000001100000000000000100000000;
		10'd152: 32'b01000101011000010000000000000000;
		10'd153: 32'b00100000000000100000000000000000;
		10'd154: 32'b00100000110000010000000000000000;
		10'd155: 32'b00000000000100000010000010000000;
		10'd156: 32'b00000000010100100000000000000000;
		10'd157: 32'b00010000000000000010000010001010;
		10'd158: 32'b11100001000000000000000000000000;
		10'd159: 32'b00000000110001000000100000000001;
		10'd160: 32'b00000000100010100001100000000000;
		10'd161: 32'b00000000000000010000100010000000;
		10'd162: 32'b00100000000000000000010000000000;
		10'd163: 32'b00001001000000000000000101000000;
		10'd164: 32'b01000000000000000000100111000010;
		10'd165: 32'b00100000000000000000000000000000;
		10'd166: 32'b00010001000000000010000000001100;
		10'd167: 32'b00010000110000010000100000000010;
		10'd168: 32'b00000100100000100010000001000000;
		10'd169: 32'b00000000000000000000000000000100;
		10'd170: 32'b00000000000000000010001000000100;
		10'd171: 32'b00000001000000000000000100011000;
		10'd172: 32'b00001000000000000000100000000100;
		10'd173: 32'b00000000000011001001000010000000;
		10'd174: 32'b00000000000010000000000001000100;
		10'd175: 32'b01000100000000000000000100000010;
		10'd176: 32'b01000000000000000000000000010000;
		10'd177: 32'b00000010000000000000000110000000;
		10'd178: 32'b00000000000000000000010000000001;
		10'd179: 32'b00000000000000000000000000000000;
		10'd180: 32'b10000000000001000000001000110000;
		10'd181: 32'b00000000000010000000000010000000;
		10'd182: 32'b10000000100000010001000000010000;
		10'd183: 32'b00100000000000000001000010000000;
		10'd184: 32'b00000000100100000000000001000100;
		10'd185: 32'b00000000101000000000000000010000;
		10'd186: 32'b00000000000000000000000110000100;
		10'd187: 32'b00000000000010000000000000100000;
		10'd188: 32'b00010000110100110001010000010001;
		10'd189: 32'b00010000000000000000001000100000;
		10'd190: 32'b00000100000001000000110100000000;
		10'd191: 32'b01000000000100000001000010000000;
		10'd192: 32'b00000001001000001000000000000000;
		10'd193: 32'b00000000001000000101001001000000;
		10'd194: 32'b00000000000000000001001000000000;
		10'd195: 32'b00000000101000000000100000000000;
		10'd196: 32'b00000000000000000000100000001000;
		10'd197: 32'b00000000000000000000000001010000;
		10'd198: 32'b00000100000010001000000000000100;
		10'd199: 32'b00000000010100000000000000000001;
		10'd200: 32'b00000000000000100100010000000000;
		10'd201: 32'b00000000000000001000000110000000;
		10'd202: 32'b00000000000000000010000000000001;
		10'd203: 32'b01000000000000000000000000010000;
		10'd204: 32'b00000000100110001000000000000000;
		10'd205: 32'b01100010000000000100000000000000;
		10'd206: 32'b00100000000001000000000000100001;
		10'd207: 32'b00000001000000100000000000001000;
		10'd208: 32'b01100000000001001000000000000000;
		10'd209: 32'b00000000000000000000110000000000;
		10'd210: 32'b00000000000100010010100010100000;
		10'd211: 32'b00010000010000100000000001000100;
		10'd212: 32'b00000001101000000000000010000010;
		10'd213: 32'b00000000000000000010000000000001;
		10'd214: 32'b00000001000001000000010000001000;
		10'd215: 32'b00000000001000000000000000000000;
		10'd216: 32'b00100100001000000011000000000100;
		10'd217: 32'b00100110000100100010000000000000;
		10'd218: 32'b00000000000010000000000000000000;
		10'd219: 32'b10000100000000000001000000001101;
		10'd220: 32'b00000000100000010000000000000000;
		10'd221: 32'b01100000011000001000000100001000;
		10'd222: 32'b10000000001001000010000000000000;
		10'd223: 32'b00010001001000000000000000000001;
		10'd224: 32'b00000100000000000000000000000000;
		10'd225: 32'b00000101000100000000100000000010;
		10'd226: 32'b00000000000111000100000010000000;
		10'd227: 32'b00000100000001001010001100000000;
		10'd228: 32'b10000000000000000000100000000000;
		10'd229: 32'b10000010000000000100000100001000;
		10'd230: 32'b00010000101000000000001010010000;
		10'd231: 32'b00000010000100100000000001000010;
		10'd232: 32'b00100000000000000000000000100000;
		10'd233: 32'b00000000100000010000010000100100;
		10'd234: 32'b00100000000000000011000010000000;
		10'd235: 32'b00000100000100000000000000000000;
		10'd236: 32'b00010000001000000000000000001000;
		10'd237: 32'b00000001010000000000000001000000;
		10'd238: 32'b10100000100100000100001010001000;
		10'd239: 32'b00000101101000000000100000000000;
		10'd240: 32'b00000000000000010000000100000000;
		10'd241: 32'b00000000000000000000010000100000;
		10'd242: 32'b10000000000000001010100110000000;
		10'd243: 32'b00000100000000000000100000000011;
		10'd244: 32'b00000000000000010010001000010001;
		10'd245: 32'b10000000000100000001000100000000;
		10'd246: 32'b00111000000000000000100000001000;
		10'd247: 32'b10000000100000000001000000011000;
		10'd248: 32'b00000000001000000000000100101000;
		10'd249: 32'b00000000000000000010000010000000;
		10'd250: 32'b00000000000000110000000000000000;
		10'd251: 32'b00000100000000110000000000000000;
		10'd252: 32'b00000000000000000000000000000001;
		10'd253: 32'b00000000000000000000000100000000;
		10'd254: 32'b01000001000000000000010001000000;
		10'd255: 32'b00000000000101000010000101000000;
		10'd256: 32'b10001000000000000010010010001100;
		10'd257: 32'b10000000000000000100010000000010;
		10'd258: 32'b00000000100000100010000000000000;
		10'd259: 32'b01000010000000000010000100000000;
		10'd260: 32'b00001000000000000001010000000101;
		10'd261: 32'b00010000010000000000110000000000;
		10'd262: 32'b00000001000000000000011000010000;
		10'd263: 32'b00101001101000000000001001001100;
		10'd264: 32'b00100000000000000000010000000000;
		10'd265: 32'b00001000000000000001000000000010;
		10'd266: 32'b00000000010000000000000000000000;
		10'd267: 32'b00000000000001000010000100000010;
		10'd268: 32'b10000000000100000100000000000000;
		10'd269: 32'b00000000000000100000000000100001;
		10'd270: 32'b00000000001100000000000000101001;
		10'd271: 32'b00000010000100000000100000000000;
		10'd272: 32'b00000000010010000100000000001000;
		10'd273: 32'b00000000000010000100000000000000;
		10'd274: 32'b00000000000100101000010000000000;
		10'd275: 32'b00010000000001001100100000100010;
		10'd276: 32'b10100101001000000000000000010000;
		10'd277: 32'b00000000000001101000000000000000;
		10'd278: 32'b00000100000000000101000000000000;
		10'd279: 32'b00000000001010100000011100010000;
		10'd280: 32'b00000001000000010000000100000001;
		10'd281: 32'b10000111000000000000000000000000;
		10'd282: 32'b10000000000000000000000100000000;
		10'd283: 32'b00000000001010010010001000000100;
		10'd284: 32'b00000000000000000000000000000000;
		10'd285: 32'b00001000000011000000000101011000;
		10'd286: 32'b10000000010000000000100010000000;
		10'd287: 32'b00000001000000000000000000000000;
		10'd288: 32'b00011000001000000000000000000001;
		10'd289: 32'b00000000100000000000000000000000;
		10'd290: 32'b01100000000100000010010000000010;
		10'd291: 32'b00000000100100000010000010000000;
		10'd292: 32'b00000000000100100000010000000010;
		10'd293: 32'b00001000000000000000000000000000;
		10'd294: 32'b00000000000100100000001001100100;
		10'd295: 32'b00100000000000000001010000000000;
		10'd296: 32'b00000100000000000000000010000110;
		10'd297: 32'b00010000010000100000000000000000;
		10'd298: 32'b10000000000010001001000000000100;
		10'd299: 32'b00000000000001000000000000000000;
		10'd300: 32'b00000000000010000000000000000000;
		10'd301: 32'b00000000000001000000100100000000;
		10'd302: 32'b01000000000000000000000010100000;
		10'd303: 32'b00000100010011000000000000000000;
		10'd304: 32'b00000000000010001001000000000100;
		10'd305: 32'b00000000000000001000000010000000;
		10'd306: 32'b00000000000000010000000000001000;
		10'd307: 32'b00100000100000000100000100000110;
		10'd308: 32'b00000000001000000000000000000100;
		10'd309: 32'b00000100010100000000000000000000;
		10'd310: 32'b00100000010001000000001000000000;
		10'd311: 32'b00100000001001000000000100100000;
		10'd312: 32'b01000000000000000100010000000000;
		10'd313: 32'b00000000000001000000000001000000;
		10'd314: 32'b10000000010000001000100000000000;
		10'd315: 32'b00000000000000000100000000000100;
		10'd316: 32'b00100000000100000001000000000000;
		10'd317: 32'b01000000100000000001000010000000;
		10'd318: 32'b00000000000000010000010000000000;
		10'd319: 32'b00000010000000000000000010000001;
		10'd320: 32'b01000001001000000000000000000000;
		10'd321: 32'b00000001000000100000000100000000;
		10'd322: 32'b00001000000010100000000000000000;
		10'd323: 32'b10000010000000000010000000000000;
		10'd324: 32'b00000000001000100000000000000000;
		10'd325: 32'b00000000000010000000000000000100;
		10'd326: 32'b10000000001010000110010000000000;
		10'd327: 32'b10000100000010000000001010100001;
		10'd328: 32'b00000000000001001000010100000100;
		10'd329: 32'b00000110001100000000000000011000;
		10'd330: 32'b00000000010000010000000101000100;
		10'd331: 32'b00000000101000001000101001000001;
		10'd332: 32'b00000000101000010000001001000010;
		10'd333: 32'b00100001000000000000000001001010;
		10'd334: 32'b00110000000001000000000000000001;
		10'd335: 32'b00000001010000000000000001000000;
		10'd336: 32'b00000000000000000000100100000000;
		10'd337: 32'b00001100000000000000010000001000;
		10'd338: 32'b00001000000000000000000000000100;
		10'd339: 32'b00000001000110010001001000000010;
		10'd340: 32'b00000001100000000010000100000000;
		10'd341: 32'b00010000000000000010000000001000;
		10'd342: 32'b11000101000000000010110000100011;
		10'd343: 32'b11000000100000000010000000000000;
		10'd344: 32'b10110010000100000000000000100000;
		10'd345: 32'b00000000000001000000000000000000;
		10'd346: 32'b00100000000000000000000000000000;
		10'd347: 32'b00000000000010001000001000000001;
		10'd348: 32'b00000000010010000100000100000000;
		10'd349: 32'b00000000000010100000000000000111;
		10'd350: 32'b00000000011000000000000000000100;
		10'd351: 32'b00000000000001000000000000000000;
		10'd352: 32'b00000011000000000000000000100000;
		10'd353: 32'b11000001110000000000000100001000;
		10'd354: 32'b00100000000000000000100000100100;
		10'd355: 32'b00101010000000000000101000000001;
		10'd356: 32'b00010000001000010000000010000000;
		10'd357: 32'b00000000000000000000000010000000;
		10'd358: 32'b00000100000001000010001000111001;
		10'd359: 32'b01000000000000000001000010001000;
		10'd360: 32'b00000000000000101000010010000000;
		10'd361: 32'b00000000000000001000000010000000;
		10'd362: 32'b00000100000000000000010000000000;
		10'd363: 32'b00010000001100000000010000100000;
		10'd364: 32'b00000000000000000000000000000000;
		10'd365: 32'b00000000101000100100000000100110;
		10'd366: 32'b00000010000011001000000000000000;
		10'd367: 32'b00100000000000000000000010000000;
		10'd368: 32'b01000000000000000000000000000000;
		10'd369: 32'b00000001000000000001000000000000;
		10'd370: 32'b00000000000000001000001100000000;
		10'd371: 32'b00100000000010000000000000100001;
		10'd372: 32'b01000100010100000001000000100000;
		10'd373: 32'b01000001000001000000110000000000;
		10'd374: 32'b10000000000000000001000101000110;
		10'd375: 32'b00000000000000000101010000100000;
		10'd376: 32'b00000100000000000100000000000010;
		10'd377: 32'b00010100100000000000000000000000;
		10'd378: 32'b00001000000000000000100001000000;
		10'd379: 32'b00000000010010000000000000000100;
		10'd380: 32'b00000000001010000000010001000000;
		10'd381: 32'b00000100000000010000000000010000;
		10'd382: 32'b00010000000100000010001010010000;
		10'd383: 32'b00010000000001000001000100100000;
		10'd384: 32'b00011000010000010000001000000100;
		10'd385: 32'b00000000000000100010000000010000;
		10'd386: 32'b00000100000010000101000000001000;
		10'd387: 32'b00001000000000001010010100110001;
		10'd388: 32'b00000010010000100000010000000000;
		10'd389: 32'b10100000100010000010010100101000;
		10'd390: 32'b00000000000000000000000000000000;
		10'd391: 32'b00001000000000000001100010000000;
		10'd392: 32'b00100010100000000000000100000000;
		10'd393: 32'b01000001000000000000000000000000;
		10'd394: 32'b00000000010000000100000010001010;
		10'd395: 32'b00100011000000000000110000001000;
		10'd396: 32'b00000100000000000000000000000000;
		10'd397: 32'b00100000000000000101000100000000;
		10'd398: 32'b00000000110010000100001000000010;
		10'd399: 32'b01010000000000010000000000000001;
		10'd400: 32'b00000100000000000110010000000010;
		10'd401: 32'b01000010010000000000100000001001;
		10'd402: 32'b00000000000100001000000000110000;
		10'd403: 32'b01000010000000000000000000000000;
		10'd404: 32'b00000000000000000000000000010100;
		10'd405: 32'b00000100000110000010010000000000;
		10'd406: 32'b00000000000000000010000000000000;
		10'd407: 32'b00000000000000110001000010000000;
		10'd408: 32'b00000100000000000100000010100100;
		10'd409: 32'b00100000100110110000000100000100;
		10'd410: 32'b00001000000000000000100010000000;
		10'd411: 32'b00000000000000000000000000000000;
		10'd412: 32'b00010100011000001001000001000000;
		10'd413: 32'b00001010000100000000000000000000;
		10'd414: 32'b00000000000000000000100100000000;
		10'd415: 32'b00010100000000000100001000000000;
		10'd416: 32'b00000000000100100000001000000000;
		10'd417: 32'b00000010010000000010000000000000;
		10'd418: 32'b00001000000011000000000010000000;
		10'd419: 32'b10000010000000000010000000000000;
		10'd420: 32'b01010000001001100000010000100110;
		10'd421: 32'b00000000000000100010010001000010;
		10'd422: 32'b00000000100000000001000000010010;
		10'd423: 32'b00001000001000000000000010010000;
		10'd424: 32'b00000000000001010000000000010100;
		10'd425: 32'b10000000000000000000000100000000;
		10'd426: 32'b00100100000001010011001100000000;
		10'd427: 32'b00000000000001010000000000000000;
		10'd428: 32'b00010000000000000000100000000000;
		10'd429: 32'b00010001000000000000000000000000;
		10'd430: 32'b00000100100010000001000000000101;
		10'd431: 32'b01000001001000000001000100000000;
		10'd432: 32'b10000010000000000100001000000000;
		10'd433: 32'b00100100000000000000000010000010;
		10'd434: 32'b01000000000000000100001000000100;
		10'd435: 32'b10000000000001000000001000000000;
		10'd436: 32'b00000000001000000000000000000000;
		10'd437: 32'b00000000000100000011000000000000;
		10'd438: 32'b10000010010000000000100000000000;
		10'd439: 32'b00000000001000010000000010001000;
		10'd440: 32'b10000000000101000000000000010010;
		10'd441: 32'b00001000000000000000101000000010;
		10'd442: 32'b00001000000000000000001000000000;
		10'd443: 32'b10000000000010000000110000000000;
		10'd444: 32'b00000000000010000000010000000000;
		10'd445: 32'b00000001000000000000000000000000;
		10'd446: 32'b00000000000100000011000101000000;
		10'd447: 32'b00000000001100000000100000100100;
		10'd448: 32'b00000000001000011010100000000100;
		10'd449: 32'b00010000000000010110100000000000;
		10'd450: 32'b00000000000000000000101000001000;
		10'd451: 32'b00000001100010001010001000100000;
		10'd452: 32'b10000000000000000001000001010010;
		10'd453: 32'b00000000010000000000000010000000;
		10'd454: 32'b00000000100000001011101000000010;
		10'd455: 32'b00000010000000000000100000100000;
		10'd456: 32'b00000000000100000000100000000000;
		10'd457: 32'b01000010000001000000000100101001;
		10'd458: 32'b00000000000000001000100010010000;
		10'd459: 32'b00000000100000000010001010000000;
		10'd460: 32'b10000000000000010000000000000000;
		10'd461: 32'b01000000000000000010000001000000;
		10'd462: 32'b00010000000000000001100000010000;
		10'd463: 32'b00000000000000000000000000000000;
		10'd464: 32'b00100000000010000000000000000000;
		10'd465: 32'b00000000000000001000000000011000;
		10'd466: 32'b00000010110001000000000010010010;
		10'd467: 32'b00100000000000001000000001000100;
		10'd468: 32'b00000000000000000000000000000000;
		10'd469: 32'b00000100000010000100000000000000;
		10'd470: 32'b00000001000000000000000100000011;
		10'd471: 32'b00000100000000100000010100000000;
		10'd472: 32'b01001100000000000000010000000000;
		10'd473: 32'b00100001000000000000100000000000;
		10'd474: 32'b00011000000000000010010000000000;
		10'd475: 32'b00000000000000001100001000100000;
		10'd476: 32'b00000010010000000100000001010000;
		10'd477: 32'b00000001000000000000000000000000;
		10'd478: 32'b00000001010000000000000000100000;
		10'd479: 32'b00000010000000000000000000000000;
		10'd480: 32'b00000000001000000000000000000000;
		10'd481: 32'b10001010000000000000101110000000;
		10'd482: 32'b00000000010000010010000001000000;
		10'd483: 32'b00010000000001000000000010010001;
		10'd484: 32'b00000000100000001000100000000100;
		10'd485: 32'b00000000000000100000000000000000;
		10'd486: 32'b00000000000100000000000000000100;
		10'd487: 32'b00010001001000000000001000100001;
		10'd488: 32'b00000000110000000000010100100000;
		10'd489: 32'b00000000000000100000000000000000;
		10'd490: 32'b00000000010000000000000000000010;
		10'd491: 32'b00101000100000001000010100000000;
		10'd492: 32'b00000000001000000000000000000000;
		10'd493: 32'b00000000000010000000000000010100;
		10'd494: 32'b00000000100000000000000000000011;
		10'd495: 32'b00000100000001000000000000010001;
		10'd496: 32'b00000000001000100000000000000010;
		10'd497: 32'b00000000000000000000001000010000;
		10'd498: 32'b00111000000000000001000000000001;
		10'd499: 32'b00000000010000000000100000000000;
		10'd500: 32'b00010000000000000101000001000000;
		10'd501: 32'b00000010100010101000000000001000;
		10'd502: 32'b00000000001000000000100000001100;
		10'd503: 32'b00000000000100000000100000101100;
		10'd504: 32'b00000001000000000000001111000010;
		10'd505: 32'b00000001000000100000100000000010;
		10'd506: 32'b00000011000000000000000110000000;
		10'd507: 32'b01001000000000000000000000000010;
		10'd508: 32'b00000100000010000000100100000000;
		10'd509: 32'b10000000000000001001000000000001;
		10'd510: 32'b00101010000100100100000100100100;
		10'd511: 32'b01100000000000000000001001000000;
		10'd512: 32'b00000001000000100000000000000000;
		10'd513: 32'b00000000000001010010000000000000;
		10'd514: 32'b00000001000001000000000000011000;
		10'd515: 32'b10100001000000000000010000001100;
		10'd516: 32'b00010000100100010000000000000010;
		10'd517: 32'b01100000000000000000001000000010;
		10'd518: 32'b00000000000000100000100000000000;
		10'd519: 32'b00010000000000000000000000000100;
		10'd520: 32'b00100000000001000000001000001000;
		10'd521: 32'b00100000001011000000000001010000;
		10'd522: 32'b10000001000100001000000000100010;
		10'd523: 32'b00000000000000000000101001000000;
		10'd524: 32'b00010010000001000010000000010000;
		10'd525: 32'b01000000001000010010100000010001;
		10'd526: 32'b00000000000000000100000000000000;
		10'd527: 32'b00000000000000000000000000000000;
		10'd528: 32'b01010010010000100000000011110010;
		10'd529: 32'b11000000000000000010000000011000;
		10'd530: 32'b10000000000000000000000000000000;
		10'd531: 32'b00000000000010000000001000000010;
		10'd532: 32'b00000100000000000001000110000000;
		10'd533: 32'b00011000000000110010010000000010;
		10'd534: 32'b00100000000100000000000000000000;
		10'd535: 32'b00000000000000001010000000000000;
		10'd536: 32'b00010000010000001001000000000100;
		10'd537: 32'b00000000010000000000000000000000;
		10'd538: 32'b00000110000000000000010000110000;
		10'd539: 32'b00000000000000000000000000000100;
		10'd540: 32'b00000000001000000000001010000000;
		10'd541: 32'b10010000000001000000000000000000;
		10'd542: 32'b00001000001000000000010000001000;
		10'd543: 32'b00000000100000001000001000000000;
		10'd544: 32'b00000000000100000110000000010000;
		10'd545: 32'b00000000000000000010000000100000;
		10'd546: 32'b00100001000000000000000000000100;
		10'd547: 32'b00010000010001000000100000000000;
		10'd548: 32'b00000000000100000010000000000100;
		10'd549: 32'b00000001000000000011110000000010;
		10'd550: 32'b00000000000000000001001000000100;
		10'd551: 32'b00000010000010000000000000000000;
		10'd552: 32'b10000001010000000000000110000000;
		10'd553: 32'b00000000010010010000100000001000;
		10'd554: 32'b11100000000010001000000100100000;
		10'd555: 32'b00000000000000010000010000000100;
		10'd556: 32'b00000110000100000100000010000000;
		10'd557: 32'b00000010000000000000100000010001;
		10'd558: 32'b10000000000000000000010000000000;
		10'd559: 32'b00011000000000000010000000010000;
		10'd560: 32'b01000010000100100000000001010000;
		10'd561: 32'b00000001101000001000000101001000;
		10'd562: 32'b00001000000000011000000000000000;
		10'd563: 32'b00000000001000110000100000000000;
		10'd564: 32'b00000000101000100000000000000000;
		10'd565: 32'b00000110000000000001000001001000;
		10'd566: 32'b00000000000000000000100000010000;
		10'd567: 32'b00000001000000000000000000010100;
		10'd568: 32'b00100010000001010000000111000000;
		10'd569: 32'b10010000010010001001000000000000;
		10'd570: 32'b00000000010000000000110000000100;
		10'd571: 32'b10000000001100000000000010000000;
		10'd572: 32'b00100001000010000001000000100000;
		10'd573: 32'b00000000000000000010000100001000;
		10'd574: 32'b01001000100000000101010000000000;
	endcase;
	return out;
endfunction
function Bit#(32) get_output_page1(UInt#(10) counter);
	Bit#(32) out = case(counter)
		10'd0: 32'b00000100100000000000000000000000;
		10'd1: 32'b00010000000100000000000000000100;
		10'd2: 32'b00000000001000000000000000100010;
		10'd3: 32'b00000001000000100000000000010000;
		10'd4: 32'b00000100000000000000000000100000;
		10'd5: 32'b10000000000000000000000000010000;
		10'd6: 32'b00000000000000000100000100010010;
		10'd7: 32'b00000000000000010000000100000010;
		10'd8: 32'b00000000000000000010000100000010;
		10'd9: 32'b00000100000001010000010000000101;
		10'd10: 32'b00000001000000010000000000000110;
		10'd11: 32'b00000001000000000000000000010010;
		10'd12: 32'b00000000000100000000000001000000;
		10'd13: 32'b00000000001000100000000000100000;
		10'd14: 32'b00000000000000000000010000100000;
		10'd15: 32'b01000000000000000001000000000000;
		10'd16: 32'b00010000000000010001000000000010;
		10'd17: 32'b00000000000000100100000000000110;
		10'd18: 32'b00000000000000010000001000000001;
		10'd19: 32'b00000000000000000101000000000110;
		10'd20: 32'b00000000000000000000000000010011;
		10'd21: 32'b00000000000000010000000000001100;
		10'd22: 32'b00000000000100010000000100010000;
		10'd23: 32'b00100000000000000000000000001000;
		10'd24: 32'b01000000000000000100000000000010;
		10'd25: 32'b00000000000000000010000000000000;
		10'd26: 32'b00000000000100000000000000010000;
		10'd27: 32'b00000000100000000000000100000010;
		10'd28: 32'b00000011000000000000000000000100;
		10'd29: 32'b00010000000000100001000000000000;
		10'd30: 32'b00010000000000000000000000000110;
		10'd31: 32'b10000000000000001000010000000000;
		10'd32: 32'b00000000010000001000000000000000;
		10'd33: 32'b00000100010000000000000001000000;
		10'd34: 32'b00000000000000000100000000001010;
		10'd35: 32'b00000001000100000000000000000100;
		10'd36: 32'b01000000010000000000000001000010;
		10'd37: 32'b00000000011000000000000000000000;
		10'd38: 32'b00010000000000100001000000000100;
		10'd39: 32'b00100000000010000000000000000000;
		10'd40: 32'b00001000000000010000000000000010;
		10'd41: 32'b00000000000000110000000000000110;
		10'd42: 32'b00000000000100100000000000000100;
		10'd43: 32'b00000000000000000010000000100000;
		10'd44: 32'b00000000000000000000000100010001;
		10'd45: 32'b00000001000000000000001000000000;
		10'd46: 32'b00000000010000000010000000000000;
		10'd47: 32'b01000000000000000000000000100000;
		10'd48: 32'b00000000000100000000000100010000;
		10'd49: 32'b00000000000001000010000000000000;
		10'd50: 32'b01010000000000100000000000000010;
		10'd51: 32'b00000000000000000100000000000001;
		10'd52: 32'b10000000000000001000010000000000;
		10'd53: 32'b00000001000000000000000000000110;
		10'd54: 32'b01010000000000000000000000000010;
		10'd55: 32'b00001000000000000001100000000000;
		10'd56: 32'b00000000000100000000000000010101;
		10'd57: 32'b00000000000000010000000100000001;
		10'd58: 32'b00000000000000010000000001000000;
		10'd59: 32'b00000000000000000000000000000110;
		10'd60: 32'b00000000000000000000000100000110;
		10'd61: 32'b00000000100001000000000010000000;
		10'd62: 32'b00000010000000010000000000000000;
		10'd63: 32'b11100011000010011010100110001000;
		10'd64: 32'b11101001010101101000010000000000;
		10'd65: 32'b00000000000010101000000001001011;
		10'd66: 32'b01101101010001001000000101000100;
		10'd67: 32'b10000000001100110110000101000000;
		10'd68: 32'b00100001001000000000000010000000;
		10'd69: 32'b01010101100000000100100000100000;
		10'd70: 32'b00100110000000011001000100101010;
		10'd71: 32'b00110100000000010101000000001001;
		10'd72: 32'b00000100100110011000110000100011;
		10'd73: 32'b01000000000001000000000100001000;
		10'd74: 32'b01100000000001100000000000001000;
		10'd75: 32'b10000100000000000000001110000000;
		10'd76: 32'b00001100000000010100000010001000;
		10'd77: 32'b10000001000000000000001101010000;
		10'd78: 32'b00100001001101101011001010101100;
		10'd79: 32'b00100000010000001010111101010000;
		10'd80: 32'b00000100000000001000010000001001;
		10'd81: 32'b00000100110000000000100001000000;
		10'd82: 32'b00000001010100000010001000000100;
		10'd83: 32'b00000010110000000000001000110010;
		10'd84: 32'b00000000000000100101010101000000;
		10'd85: 32'b10001000010010000001010001111000;
		10'd86: 32'b00000000000000100000001000000010;
		10'd87: 32'b00000100000001010010000011000001;
		10'd88: 32'b00011101101001110100100101010000;
		10'd89: 32'b01000110000111000010001010100001;
		10'd90: 32'b10010000000011000010001100000000;
		10'd91: 32'b00000000000010000010010000000000;
		10'd92: 32'b00000100110000000000000001001000;
		10'd93: 32'b00010000000101001000010000110010;
		10'd94: 32'b01000010101000000001110100010010;
		10'd95: 32'b01100100000100000010010011000000;
		10'd96: 32'b00000000000100010000000000000000;
		10'd97: 32'b10001010000101011000010010001000;
		10'd98: 32'b00110000101001010101001000000000;
		10'd99: 32'b00000100000000000010010000000100;
		10'd100: 32'b01001000100001010100000000000000;
		10'd101: 32'b01000000000001100000011000001011;
		10'd102: 32'b00101100000000011000000001000001;
		10'd103: 32'b00001010100000000011000000000101;
		10'd104: 32'b00000010110101000110000100000000;
		10'd105: 32'b00001110010101001000000000010000;
		10'd106: 32'b00000010000000100110100010000011;
		10'd107: 32'b00101001100000111000001100000100;
		10'd108: 32'b00000110010100011010001000001000;
		10'd109: 32'b00001010001000101100000100000001;
		10'd110: 32'b01000000000000000000001001101000;
		10'd111: 32'b00111100100001100000010000100000;
		10'd112: 32'b10110100000001000100001100000101;
		10'd113: 32'b00000100000100000111100000010000;
		10'd114: 32'b10100011000001100000110001100000;
		10'd115: 32'b00100100000010101000000001000000;
		10'd116: 32'b11100010111000001010010000010001;
		10'd117: 32'b00011010000000100110001001000100;
		10'd118: 32'b00011000000010000000100000100010;
		10'd119: 32'b00100000010000100001000001000000;
		10'd120: 32'b00010100000000001001000011010010;
		10'd121: 32'b01100110000000100000000000011111;
		10'd122: 32'b00000000010100000001010001100001;
		10'd123: 32'b00100000000000000001101010010010;
		10'd124: 32'b00001000010001010000100100000100;
		10'd125: 32'b00000010001010000100000100000000;
		10'd126: 32'b11001011000100010100100100100011;
		10'd127: 32'b00101001000010000110000100000001;
		10'd128: 32'b00110000100100011000000000000010;
		10'd129: 32'b00000000000011000011000010011100;
		10'd130: 32'b00000010001110101000000011100011;
		10'd131: 32'b01001101000010000100000001110001;
		10'd132: 32'b00011000100100001000100010000010;
		10'd133: 32'b00100000101010000001000011001000;
		10'd134: 32'b01011010011011000001100000010110;
		10'd135: 32'b10101001001000001000000110101000;
		10'd136: 32'b01011001000000010000000000100000;
		10'd137: 32'b10000100010000101000100000001101;
		10'd138: 32'b10110001110001000000100010000001;
		10'd139: 32'b10000000100000000000110000000010;
		10'd140: 32'b00101000000010000000001100100000;
		10'd141: 32'b00010111000000111000111100001100;
		10'd142: 32'b01000010100011000001001000000000;
		10'd143: 32'b00010100000000010100000000010000;
		10'd144: 32'b01000000110011001000000010001010;
		10'd145: 32'b00000100000100100001110000000000;
		10'd146: 32'b01100100010010101100100010000000;
		10'd147: 32'b00100100001010001100001000000001;
		10'd148: 32'b00101000000100010100000011000101;
		10'd149: 32'b00100010000000000101001001000000;
		10'd150: 32'b10100000101000000100100011101000;
		10'd151: 32'b00000001100000000010000100000000;
		10'd152: 32'b01000101011000010000010000000000;
		10'd153: 32'b00100000000001101010000000000010;
		10'd154: 32'b00100000110001010000000000110000;
		10'd155: 32'b00000001000100000010000110001000;
		10'd156: 32'b01111011010100110100000000000000;
		10'd157: 32'b00110000000000000010000010001010;
		10'd158: 32'b11100001110000000100000000001100;
		10'd159: 32'b00000000110001000000100000101001;
		10'd160: 32'b00100010100110100101100001000000;
		10'd161: 32'b10000000100000010000100010001010;
		10'd162: 32'b00110100100100000000011000000000;
		10'd163: 32'b00001111000001000010000101000010;
		10'd164: 32'b01000000111101000000101111101010;
		10'd165: 32'b00100000100100000000110000000001;
		10'd166: 32'b01010001100000000010000000001100;
		10'd167: 32'b00010110110000010001100100000010;
		10'd168: 32'b01000100110000100010000101000110;
		10'd169: 32'b00011000010011000000000010000100;
		10'd170: 32'b00000000100010000010011000010100;
		10'd171: 32'b00000001000000000100010100011010;
		10'd172: 32'b00101100000000001000110000010100;
		10'd173: 32'b00000000001011111001010010000000;
		10'd174: 32'b00000000100011000000110001000100;
		10'd175: 32'b01100101000000000000001100100010;
		10'd176: 32'b01000000000000100010111000010000;
		10'd177: 32'b10000010000000000000001110100001;
		10'd178: 32'b00000000000000000000010001011001;
		10'd179: 32'b00000100000000000000000001011000;
		10'd180: 32'b11000010001001000101001000111000;
		10'd181: 32'b00001010001110000001100110000000;
		10'd182: 32'b10000010100000010001000000110000;
		10'd183: 32'b01110000000000001001000010100010;
		10'd184: 32'b00000110101100010000110001101100;
		10'd185: 32'b00000000101000000000000100010000;
		10'd186: 32'b00100000000001001000100110000100;
		10'd187: 32'b01000010000010010000001000100000;
		10'd188: 32'b00010000110101111001010000010101;
		10'd189: 32'b00010000000000001000011100100010;
		10'd190: 32'b01100100100101000000110100000000;
		10'd191: 32'b01000100010100100001001110010001;
		10'd192: 32'b00000001001000001100000010000101;
		10'd193: 32'b00000000011100000101001001000000;
		10'd194: 32'b00000000000000000001101000100010;
		10'd195: 32'b00000000101000010010111000000011;
		10'd196: 32'b01000000010000000000110000011000;
		10'd197: 32'b00101000000110001000000001010000;
		10'd198: 32'b00110100000010001000000000001100;
		10'd199: 32'b00000000010100010000000001000001;
		10'd200: 32'b00000000000100100100010010000000;
		10'd201: 32'b01100000100000001000000110011000;
		10'd202: 32'b00110000010100000110000000000001;
		10'd203: 32'b01000000010000010001000000010000;
		10'd204: 32'b01100000100110011010000001010000;
		10'd205: 32'b01110010100000000101000000000000;
		10'd206: 32'b00100100000001000100000001100001;
		10'd207: 32'b01000001000010101000000110001000;
		10'd208: 32'b01100010000001001010000001000010;
		10'd209: 32'b00000101000000000000110010100000;
		10'd210: 32'b00000000100110010010110010100000;
		10'd211: 32'b00010010110000111000001101000110;
		10'd212: 32'b00000011101100010000101010000010;
		10'd213: 32'b00001000000000000010000000001001;
		10'd214: 32'b00000001001001000000010000101001;
		10'd215: 32'b00000000011000011000000000000000;
		10'd216: 32'b10100101001000000011000010000100;
		10'd217: 32'b00100110000100101010001010000000;
		10'd218: 32'b00010000001010010000000000000000;
		10'd219: 32'b10000100110110101011000000011101;
		10'd220: 32'b00000000110000010000000101000000;
		10'd221: 32'b01111000011001001000000110001100;
		10'd222: 32'b10000000001001000010000000000110;
		10'd223: 32'b00010011001000000000000000000001;
		10'd224: 32'b00000100010000000000001000000000;
		10'd225: 32'b01001101000101101000100110000010;
		10'd226: 32'b00000001000111100101000110000100;
		10'd227: 32'b00000101000101111010001110000000;
		10'd228: 32'b10000010000000001000100000010000;
		10'd229: 32'b10100010000000010100100100001000;
		10'd230: 32'b01010000101000000100001010010000;
		10'd231: 32'b00000010000100101000000001000010;
		10'd232: 32'b00100000001100000011001000100010;
		10'd233: 32'b00000000100000010000011100101110;
		10'd234: 32'b01100100000000000111000010000000;
		10'd235: 32'b00000100000100000000000000000000;
		10'd236: 32'b00110100101000000000000000001000;
		10'd237: 32'b10001001010100000000100101011100;
		10'd238: 32'b10100000100110000100001010001000;
		10'd239: 32'b00000101101000100000100110010000;
		10'd240: 32'b00000000000000010000100100000010;
		10'd241: 32'b00110000100000000000010011110100;
		10'd242: 32'b10001100000001001010100110000000;
		10'd243: 32'b00000100000010000100100100000011;
		10'd244: 32'b00000000000100010110001010010001;
		10'd245: 32'b10000000101100010001100110100100;
		10'd246: 32'b00111100100000000011100010001000;
		10'd247: 32'b10000011100000000001000010011010;
		10'd248: 32'b01000100101000000000000110101010;
		10'd249: 32'b00000000000001100010000010010000;
		10'd250: 32'b10010001100100110000000000000000;
		10'd251: 32'b00000100000000110001000010000000;
		10'd252: 32'b00000000010000000000000011001011;
		10'd253: 32'b01000000000011010000000110011000;
		10'd254: 32'b01000011001000000001010111001000;
		10'd255: 32'b00000000010111001010000101000000;
		10'd256: 32'b10001000110000000010010010011101;
		10'd257: 32'b11000000010000001110010000000010;
		10'd258: 32'b10001000100000100011000000000000;
		10'd259: 32'b01001010001000001010101101000000;
		10'd260: 32'b10001010100000000101010110001101;
		10'd261: 32'b00010100010001000000110000000000;
		10'd262: 32'b00000001010000000010011000010100;
		10'd263: 32'b00111001101100000000101001001100;
		10'd264: 32'b00110000000000000000110000010000;
		10'd265: 32'b10001000000000000001100000010011;
		10'd266: 32'b01000000010000000000000011010000;
		10'd267: 32'b00100000000001000010000100000010;
		10'd268: 32'b10001001010100000100000010001000;
		10'd269: 32'b00000000010000100111100010110111;
		10'd270: 32'b00000000001100001000100000101101;
		10'd271: 32'b00000010010100000100100100001000;
		10'd272: 32'b00001100011011000110000000001000;
		10'd273: 32'b01000100100010000100000000000010;
		10'd274: 32'b00000000010100101001010001000000;
		10'd275: 32'b01110011100001001100100100100010;
		10'd276: 32'b11100101011000001001000100010000;
		10'd277: 32'b00000010100011101000100000000010;
		10'd278: 32'b01000100010001000101000000000000;
		10'd279: 32'b10010000001010100000011100010000;
		10'd280: 32'b01000101000000010001000101000001;
		10'd281: 32'b10100111101000000000000000000001;
		10'd282: 32'b11100000000100000010001100010000;
		10'd283: 32'b00000000001010010010011010100100;
		10'd284: 32'b11001010100000001000000010000000;
		10'd285: 32'b00001000000011010000000111011000;
		10'd286: 32'b10000010110010011000100010010000;
		10'd287: 32'b00000001010100001000100000100000;
		10'd288: 32'b00011000001100001100010000000101;
		10'd289: 32'b10001000100000000000010100000000;
		10'd290: 32'b01110000001100000010010000000011;
		10'd291: 32'b00011001110100100010000010000000;
		10'd292: 32'b10100001011100101010010000000011;
		10'd293: 32'b01001010010000000001010101000000;
		10'd294: 32'b10000001000100100000001001110100;
		10'd295: 32'b00100000011010000011110010001010;
		10'd296: 32'b00010100000010100101000010100110;
		10'd297: 32'b01010000110001100000010001000000;
		10'd298: 32'b11000000000010001001000000100100;
		10'd299: 32'b00000010000001000000110000000000;
		10'd300: 32'b11000010000010000000000000000000;
		10'd301: 32'b00000100001001001101100100000000;
		10'd302: 32'b01000001110010000000000010100000;
		10'd303: 32'b10000100110011100000100000000000;
		10'd304: 32'b00010000000010001001000100000100;
		10'd305: 32'b00000011000001011100000010000000;
		10'd306: 32'b00000100000000110000001000001001;
		10'd307: 32'b01101000100001100100000100010110;
		10'd308: 32'b00000001001001000000001000000100;
		10'd309: 32'b00010101010100010010000000001000;
		10'd310: 32'b00101000010001000000101000111010;
		10'd311: 32'b00100000001001000001000100100000;
		10'd312: 32'b01000000001000000100010010000000;
		10'd313: 32'b00000000000001010000100001000000;
		10'd314: 32'b10010000010000101010100000000000;
		10'd315: 32'b00000100000001000100000010000100;
		10'd316: 32'b00110000100101000001000000000001;
		10'd317: 32'b01100001101000010011000110000000;
		10'd318: 32'b00010010011010010000010000000000;
		10'd319: 32'b00000010000000000001000110010001;
		10'd320: 32'b01001001001000010010001000000000;
		10'd321: 32'b10000001001000111000001100001100;
		10'd322: 32'b00011110000010100000000000000000;
		10'd323: 32'b10010010010000010010000000000000;
		10'd324: 32'b00010010001000100000101000000000;
		10'd325: 32'b00000000001010000000000001110100;
		10'd326: 32'b10000000111010000110010000000000;
		10'd327: 32'b10000100100010001000001010110001;
		10'd328: 32'b00000000001001011010011100000101;
		10'd329: 32'b00101110001100000000000001111000;
		10'd330: 32'b00000000010000010100010101010101;
		10'd331: 32'b00000010101000011000101001000001;
		10'd332: 32'b10100100111110011000011101000010;
		10'd333: 32'b00110001000010000000000001001011;
		10'd334: 32'b00110101010001000000000100000001;
		10'd335: 32'b00000001010000000000110001001000;
		10'd336: 32'b00000100010000000000100100100100;
		10'd337: 32'b00011101010000000000010000001000;
		10'd338: 32'b01001000001000000000010000001101;
		10'd339: 32'b10000001010110010101001000001011;
		10'd340: 32'b00000001101000000110100100001001;
		10'd341: 32'b00110000000000000011000001001000;
		10'd342: 32'b11000101001000000010110100100011;
		10'd343: 32'b11001100110110000010000000000001;
		10'd344: 32'b10110010010100110000000010100000;
		10'd345: 32'b00001000010001100010100000000011;
		10'd346: 32'b10100001001000000100000110000001;
		10'd347: 32'b11000000000010011000001000010001;
		10'd348: 32'b00000000010010001100010100100000;
		10'd349: 32'b00000000100010110000010000000111;
		10'd350: 32'b00000000011000000000000000000100;
		10'd351: 32'b11100100001001000010001010001000;
		10'd352: 32'b00100111100001010001000000110000;
		10'd353: 32'b11000001110000000010000110001000;
		10'd354: 32'b00100000110000000000110001100100;
		10'd355: 32'b00101010000000000000101000101011;
		10'd356: 32'b00010001101000010000000011000001;
		10'd357: 32'b00000000010000000001000010000001;
		10'd358: 32'b00000110100001001010001000111001;
		10'd359: 32'b11101001000000001001010110001000;
		10'd360: 32'b10000010000000101110010010000000;
		10'd361: 32'b01000010000100001000000010000000;
		10'd362: 32'b00011110000000000100010000001000;
		10'd363: 32'b10011000001100001010010100100000;
		10'd364: 32'b00000001000110001000000000000010;
		10'd365: 32'b00000000111000100110000000100110;
		10'd366: 32'b01000010000111001110000001000000;
		10'd367: 32'b00100000101011101000001010100000;
		10'd368: 32'b01010010000100100000000001000000;
		10'd369: 32'b01011001001010000001000000000000;
		10'd370: 32'b00000001000000001001001100000000;
		10'd371: 32'b00100000001010110000000110100001;
		10'd372: 32'b11001100110100000001000000100000;
		10'd373: 32'b11100001010101000100110000000001;
		10'd374: 32'b10000000000000000001001101100110;
		10'd375: 32'b10000000000000000101010000110000;
		10'd376: 32'b00000101000000000100000001001110;
		10'd377: 32'b01010100100100000000000001010101;
		10'd378: 32'b00011001000000000000101011010000;
		10'd379: 32'b01001000110010000001000000000100;
		10'd380: 32'b00011001001010000100110001000010;
		10'd381: 32'b00101100000000110010000000010011;
		10'd382: 32'b00110100000100000011001011010000;
		10'd383: 32'b10010000000001000001000100100000;
		10'd384: 32'b00011110010100011100001001000100;
		10'd385: 32'b00000100010100100010000000110000;
		10'd386: 32'b00000100000010010101000000001010;
		10'd387: 32'b00011100001000001011010100110011;
		10'd388: 32'b10000010011000100000010001000000;
		10'd389: 32'b10100001100010000010010100101000;
		10'd390: 32'b11000010001010000000000000000000;
		10'd391: 32'b01001000000000000011100011001001;
		10'd392: 32'b01100010100000100000000100000010;
		10'd393: 32'b01000011010000000010010000101110;
		10'd394: 32'b00000000011100000101001011001010;
		10'd395: 32'b01110011100010001000110000001100;
		10'd396: 32'b00100100010000010101000000000010;
		10'd397: 32'b10100100010000000101001100000000;
		10'd398: 32'b00000011110010000100001000000010;
		10'd399: 32'b01010010010000010000010000000001;
		10'd400: 32'b10000100010000000110110100100110;
		10'd401: 32'b01000010010000000000100000001001;
		10'd402: 32'b00000000010100001000000000111000;
		10'd403: 32'b01000011000000000000010000011000;
		10'd404: 32'b00000000100000100010000010010101;
		10'd405: 32'b01010100000110110010010000000000;
		10'd406: 32'b00010100010000000110001000100010;
		10'd407: 32'b00001000100100110011000110000000;
		10'd408: 32'b00010100100000000100000011100100;
		10'd409: 32'b00100100100111110100110100000100;
		10'd410: 32'b00001000000100100000100010000000;
		10'd411: 32'b01000000000000000000101000010000;
		10'd412: 32'b10110110011000101001010001001000;
		10'd413: 32'b00001011000110000000000000000000;
		10'd414: 32'b10000000000000000000110100000000;
		10'd415: 32'b00110110001000000100001000000000;
		10'd416: 32'b10000000000111100000011001010000;
		10'd417: 32'b00000010010100100010000000000000;
		10'd418: 32'b00001000001011000011000110011000;
		10'd419: 32'b10000010000000000011100100000100;
		10'd420: 32'b01010000001011100000010000110110;
		10'd421: 32'b00001000000000100010010101000010;
		10'd422: 32'b10000100101000100001100000010010;
		10'd423: 32'b00001000001000100010000010010000;
		10'd424: 32'b00100000000001010000000100010100;
		10'd425: 32'b10000000000000000000100100010100;
		10'd426: 32'b00100100000011010011001110000000;
		10'd427: 32'b10000000001101010000000010000001;
		10'd428: 32'b00110000000011010000100000000000;
		10'd429: 32'b00111001000000000000000000000100;
		10'd430: 32'b10000100101010010001011100010111;
		10'd431: 32'b11110101001000000011000100000000;
		10'd432: 32'b10000010100000000100001001000110;
		10'd433: 32'b00100101001100000010000010000010;
		10'd434: 32'b11001000001000000100001100000100;
		10'd435: 32'b10000000100001000100001000000000;
		10'd436: 32'b00000000001000000100010000000000;
		10'd437: 32'b00100000000100000011100000001000;
		10'd438: 32'b10000010110000000111111000000000;
		10'd439: 32'b10000001001010010000010010001010;
		10'd440: 32'b10001000000101100001001000010010;
		10'd441: 32'b00001001000000000000101001000110;
		10'd442: 32'b00001000000000000011011100000000;
		10'd443: 32'b10000010000010000000110000000010;
		10'd444: 32'b00000000000010100101010000000001;
		10'd445: 32'b00010001001000001000000000100010;
		10'd446: 32'b01010000000110010011010111000110;
		10'd447: 32'b00000000001100000000100000100100;
		10'd448: 32'b00010000001000011110100101000110;
		10'd449: 32'b01010000001000010111100010000101;
		10'd450: 32'b00000000000000000100101000011000;
		10'd451: 32'b00000001100010011111111000100000;
		10'd452: 32'b10100001001000000001001011010010;
		10'd453: 32'b00010000011000000000001010000000;
		10'd454: 32'b11010000100000001011101000000010;
		10'd455: 32'b00000010001000000000100000100111;
		10'd456: 32'b00001000000100000000100100000000;
		10'd457: 32'b01000010000001001000000100111001;
		10'd458: 32'b00000000000000001000100010011000;
		10'd459: 32'b00101110100000010011001010010100;
		10'd460: 32'b10000010000000110000000100000000;
		10'd461: 32'b11000000001000000010000101010000;
		10'd462: 32'b00011000000000000011100000010000;
		10'd463: 32'b00100000000000000100011000000000;
		10'd464: 32'b00100000010110001000000000000000;
		10'd465: 32'b00000000001010001000000010011000;
		10'd466: 32'b00010010110001101000000010011010;
		10'd467: 32'b00100100000010101000010001010110;
		10'd468: 32'b00000100000000001000000000001000;
		10'd469: 32'b00000100010010000100000000000000;
		10'd470: 32'b01010101011001010000000101001011;
		10'd471: 32'b00000100000000100010010100100000;
		10'd472: 32'b01011101000010100000010000010000;
		10'd473: 32'b00100001000010000010100000010001;
		10'd474: 32'b00011001100001000110110000000000;
		10'd475: 32'b00000011000100101100001000100100;
		10'd476: 32'b00000110010001000101000001110000;
		10'd477: 32'b01001001000000001010000000100000;
		10'd478: 32'b00001011010000000110001000101000;
		10'd479: 32'b00100010000000000000001010000000;
		10'd480: 32'b00000000011000000000000101000000;
		10'd481: 32'b10101110000000001000101110000000;
		10'd482: 32'b00100100010000010010000001000000;
		10'd483: 32'b01010000001001000100110010110101;
		10'd484: 32'b10100000101001001000100000000110;
		10'd485: 32'b00001000000000101000000000011000;
		10'd486: 32'b00000000000101000000010100001100;
		10'd487: 32'b10110001001100000000001000100001;
		10'd488: 32'b00100010110000000000010100100010;
		10'd489: 32'b11100001000000100000000000000000;
		10'd490: 32'b00000000110000101000000001000011;
		10'd491: 32'b00101000110000011000010100001010;
		10'd492: 32'b00001010101000100000000000000000;
		10'd493: 32'b00000000000010001000100000011100;
		10'd494: 32'b00001000100000011001010000000011;
		10'd495: 32'b00000100000001010000000100010001;
		10'd496: 32'b10000000001000100100000000100110;
		10'd497: 32'b00000000001010010000011000010100;
		10'd498: 32'b00111000101100100001000000100101;
		10'd499: 32'b00010001010011000100100000000001;
		10'd500: 32'b00010000001000001111000001100100;
		10'd501: 32'b01000010100010101000010000001000;
		10'd502: 32'b00100000001010000010101000001100;
		10'd503: 32'b01000000100100000000100000101111;
		10'd504: 32'b00000111101000001000001111000110;
		10'd505: 32'b10000001101000110001100000000011;
		10'd506: 32'b00000011011100000000000110000010;
		10'd507: 32'b01001100000000000000100000010010;
		10'd508: 32'b00001100000010000000111100000000;
		10'd509: 32'b10000000000100001001000000000001;
		10'd510: 32'b10101010001101100110000100101101;
		10'd511: 32'b01100000001000100000001001001000;
		10'd512: 32'b01000101001000100000100001000010;
		10'd513: 32'b00001001000001010010000100100010;
		10'd514: 32'b10000001000001001000001000011000;
		10'd515: 32'b11100001000000000001010010001100;
		10'd516: 32'b01011000100101010000000000000010;
		10'd517: 32'b01101001000000000000001010000010;
		10'd518: 32'b10100100000001100010100000010000;
		10'd519: 32'b00011101001000000010000000000101;
		10'd520: 32'b00110001000001000001001000001000;
		10'd521: 32'b00101100001011000000000001011000;
		10'd522: 32'b11000001100100101000010000110010;
		10'd523: 32'b00001010110000000100101001100000;
		10'd524: 32'b01011010000111000011100000010010;
		10'd525: 32'b01001000001001110110100100010011;
		10'd526: 32'b11000000000100000100000100100000;
		10'd527: 32'b00000001000010000001000000000100;
		10'd528: 32'b01010010010000100001000111111010;
		10'd529: 32'b11010000000001000110001000011010;
		10'd530: 32'b10000000000000000000000100000010;
		10'd531: 32'b10000000000010000001001000100010;
		10'd532: 32'b00001101001000000001001110000000;
		10'd533: 32'b00011000000001110010010010110011;
		10'd534: 32'b00101000001111100000000010000000;
		10'd535: 32'b00000001000000001011111000000100;
		10'd536: 32'b00010001010000001001000010001100;
		10'd537: 32'b00000010010011001000000000100000;
		10'd538: 32'b00000110001000010000110000110001;
		10'd539: 32'b00100001000110000000010000000100;
		10'd540: 32'b00100000001000000010001010100000;
		10'd541: 32'b10010000000001000110000000000001;
		10'd542: 32'b00001000001000000100110011001111;
		10'd543: 32'b01010000100000001000001000000100;
		10'd544: 32'b00000000010100000110100101110000;
		10'd545: 32'b10000010000100010010000000100001;
		10'd546: 32'b00100001010000000000001001000100;
		10'd547: 32'b00010000010011000000100000000000;
		10'd548: 32'b00000100100100000010000001000100;
		10'd549: 32'b00000101000000000011110000000010;
		10'd550: 32'b00000001010000011001001000000100;
		10'd551: 32'b00000011000010010000110000000000;
		10'd552: 32'b10101001110000101100000110000000;
		10'd553: 32'b00000000011110110010100100101000;
		10'd554: 32'b11100000000110001000000110100000;
		10'd555: 32'b00010001000000010101010000100100;
		10'd556: 32'b00000110000110000100000010000000;
		10'd557: 32'b01000010110110000000100000111001;
		10'd558: 32'b11011001000100000100010001001000;
		10'd559: 32'b01011000000000000011000000010000;
		10'd560: 32'b01000010001100100000000001010010;
		10'd561: 32'b01010001101000001000000101001000;
		10'd562: 32'b00101000000001111000100001000000;
		10'd563: 32'b00001000001010111010100010001000;
		10'd564: 32'b00000000101000100000000000000000;
		10'd565: 32'b00000111000000000001000001001101;
		10'd566: 32'b00001000001000010000100001010100;
		10'd567: 32'b00000101000000000000010000010100;
		10'd568: 32'b01110010100001010000000111000000;
		10'd569: 32'b10010011110010011001100100000000;
		10'd570: 32'b01100000011000000001110001000110;
		10'd571: 32'b10000001101101000000000010100000;
		10'd572: 32'b00100001000010000001010010110000;
		10'd573: 32'b00101000100001001010010100001000;
		10'd574: 32'b01001000100000000101110000000000;
	endcase;
	return out;
endfunction
function Bit#(32) get_output_page2(UInt#(10) counter);
	Bit#(32) out = case(counter)
		10'd0: 32'b00000100100000000100000010000000;
		10'd1: 32'b00010000000100000000000000100100;
		10'd2: 32'b00000000001000000000000001100010;
		10'd3: 32'b00000001000000100000000001010010;
		10'd4: 32'b00000100000000000100000000100000;
		10'd5: 32'b10000000000000010000000000010000;
		10'd6: 32'b01000000000000100100000100010010;
		10'd7: 32'b00000000000000010001000100000110;
		10'd8: 32'b00000100000000000010000100000010;
		10'd9: 32'b00000101000001010000010000010101;
		10'd10: 32'b00000001000000010000000000000110;
		10'd11: 32'b00010001000000000000000000010010;
		10'd12: 32'b00000000010100000000000101000000;
		10'd13: 32'b00000000001000100000000000110100;
		10'd14: 32'b00000100000100000000010000100000;
		10'd15: 32'b01000000000000000101000100000000;
		10'd16: 32'b00010000010000110001000000000010;
		10'd17: 32'b01100000000001100110000000000110;
		10'd18: 32'b00000000000000010000001010000001;
		10'd19: 32'b00000000000000010101000000000111;
		10'd20: 32'b00000000000001100000000000010011;
		10'd21: 32'b00000000001000010000000000001100;
		10'd22: 32'b00000000000100010000000100010000;
		10'd23: 32'b00100000000000000000000000101000;
		10'd24: 32'b01000000000000000100000100000010;
		10'd25: 32'b00100000001000000010000000100000;
		10'd26: 32'b00100000000100000000000000010000;
		10'd27: 32'b00000000110000100000000111000010;
		10'd28: 32'b00000011000000000001000000000100;
		10'd29: 32'b00010100000000100001000000000000;
		10'd30: 32'b00010000000000000001000100000110;
		10'd31: 32'b10000000000100001000010000000000;
		10'd32: 32'b10000000010000001001000000000000;
		10'd33: 32'b01000100010000000000001001000000;
		10'd34: 32'b00010000000000000100000000001010;
		10'd35: 32'b00000001000100000000000100000101;
		10'd36: 32'b01000000010100000000000001000010;
		10'd37: 32'b00000000011000000001000001000000;
		10'd38: 32'b00010000000000100001001000000100;
		10'd39: 32'b00100000000010000000000000000010;
		10'd40: 32'b00011000000000010000100000000010;
		10'd41: 32'b00000010000000110100000000000110;
		10'd42: 32'b01000000000100100000000000000110;
		10'd43: 32'b00000000000000000110001000100000;
		10'd44: 32'b00100000000000000000000100010001;
		10'd45: 32'b00000001000100000000001100000000;
		10'd46: 32'b00000000010000010010000001000000;
		10'd47: 32'b11000000000010000000000000100000;
		10'd48: 32'b00000000100100000000000100010000;
		10'd49: 32'b10100000000001001010000000000000;
		10'd50: 32'b01010000000000100000010000000110;
		10'd51: 32'b00000001000000000100000100000001;
		10'd52: 32'b10000100000000101000010000000000;
		10'd53: 32'b00000101000001000000010000000110;
		10'd54: 32'b01010000000001000000000000000110;
		10'd55: 32'b00001000000000000001100000001000;
		10'd56: 32'b00000000000100000000000010010101;
		10'd57: 32'b00000001000000110000000100000001;
		10'd58: 32'b00010000010000010000000001000000;
		10'd59: 32'b00000000000001100000000000000110;
		10'd60: 32'b00000000000000100001000100000110;
		10'd61: 32'b00000000100001000010000010000000;
		10'd62: 32'b00000010000000010000000000010001;
		10'd63: 32'b11110011000010011010100110001001;
		10'd64: 32'b11101111110111101000010100001000;
		10'd65: 32'b11000000010010101000000101101011;
		10'd66: 32'b11111101110001001000000101000101;
		10'd67: 32'b10000001011110110110010101000000;
		10'd68: 32'b01100011001110100100000010010000;
		10'd69: 32'b01010101100010000110100001110000;
		10'd70: 32'b10100111000000011011011100101011;
		10'd71: 32'b00110110000000010101000000001001;
		10'd72: 32'b10000101100110011000110100101011;
		10'd73: 32'b11000100001001010000010100001100;
		10'd74: 32'b11100000000101100000001000001000;
		10'd75: 32'b10000101000000110010011110000000;
		10'd76: 32'b10111100010010010101001110001001;
		10'd77: 32'b10000001000011000001001101010000;
		10'd78: 32'b11110101001101101011001110101101;
		10'd79: 32'b11101010011000001010111101110001;
		10'd80: 32'b01000100000101011000011001001001;
		10'd81: 32'b00000110111000100010110001000010;
		10'd82: 32'b00000001011100000010011000000100;
		10'd83: 32'b10000010111101000101001000110010;
		10'd84: 32'b01000110000010110111010101000001;
		10'd85: 32'b10001000011010000001010001111100;
		10'd86: 32'b01000000001110100010001000100110;
		10'd87: 32'b00100100001011010010000111000001;
		10'd88: 32'b00011101101011111110100101010000;
		10'd89: 32'b01000110000111010011001010100101;
		10'd90: 32'b10110000001011100011001110000010;
		10'd91: 32'b00100101000010000010011000000011;
		10'd92: 32'b00000111110101100000100001101011;
		10'd93: 32'b00110100010101001100011100110011;
		10'd94: 32'b01000010101001000001111100010111;
		10'd95: 32'b01100100010101010010010111001011;
		10'd96: 32'b00011000000101010100000000000001;
		10'd97: 32'b10001011000101011000110010001101;
		10'd98: 32'b00110000101011110101011100000101;
		10'd99: 32'b11000100010000010110010000000100;
		10'd100: 32'b01101010111001010100001000000000;
		10'd101: 32'b01000001010001110000011000001011;
		10'd102: 32'b00111100000000011001000101000001;
		10'd103: 32'b10101111100000000011000010000101;
		10'd104: 32'b11010010110101101110000100101100;
		10'd105: 32'b00011110011101101000010100010000;
		10'd106: 32'b00000010010110100110100010000011;
		10'd107: 32'b00101011100100111000001110000100;
		10'd108: 32'b00010111111101011010111100011000;
		10'd109: 32'b00001011111010101100000101010101;
		10'd110: 32'b01001010000010000000001001101001;
		10'd111: 32'b00111100101011110001010010101010;
		10'd112: 32'b11110100000001100110001101010111;
		10'd113: 32'b00000100000100000111100000110010;
		10'd114: 32'b10110011000101101100110001101010;
		10'd115: 32'b00100110000010111100001001100000;
		10'd116: 32'b11100010111001001010010000010001;
		10'd117: 32'b00011010000100100111001001010100;
		10'd118: 32'b11011000000110100000100010100011;
		10'd119: 32'b00111000010100100001000001010110;
		10'd120: 32'b10010100000000011001000011010010;
		10'd121: 32'b01100110000100100001000000011111;
		10'd122: 32'b10100101010100000001010001101101;
		10'd123: 32'b00101000000000000011101011010010;
		10'd124: 32'b00011000010001011000100100110100;
		10'd125: 32'b00110111011010000100000100010110;
		10'd126: 32'b11011011100100010100100110111011;
		10'd127: 32'b01111011001010001111001110010001;
		10'd128: 32'b00111000100100111100010000000010;
		10'd129: 32'b00000000001111000111001010011101;
		10'd130: 32'b00100011001110101010000011110111;
		10'd131: 32'b01001101000010000100000001110001;
		10'd132: 32'b10011000101101001010100010000010;
		10'd133: 32'b00100000101011000001000011011100;
		10'd134: 32'b11111010011011101001100001011111;
		10'd135: 32'b10111101001000001000100111101000;
		10'd136: 32'b11111101000100011000100000100000;
		10'd137: 32'b10000100010001111000100000001101;
		10'd138: 32'b10110111110111000000100110000001;
		10'd139: 32'b10001100100000000011110000100010;
		10'd140: 32'b00101010000110000000101100110000;
		10'd141: 32'b00010111010000111010111110001101;
		10'd142: 32'b11101011110011100001001100001000;
		10'd143: 32'b00110100001100010100000000010000;
		10'd144: 32'b01000000111011001000100010111010;
		10'd145: 32'b00100100000100100001110000001000;
		10'd146: 32'b11111101010010111100100010001001;
		10'd147: 32'b00100100001010001101111100010001;
		10'd148: 32'b00101000000101010110000011100111;
		10'd149: 32'b00100010000000011101011001010000;
		10'd150: 32'b10110010101010000100100011101000;
		10'd151: 32'b10000001100001000110000110001000;
		10'd152: 32'b11001101111100011000010110000000;
		10'd153: 32'b00100000000001101010000000001010;
		10'd154: 32'b01100001110001011000000000111000;
		10'd155: 32'b00000011100101000110000110011010;
		10'd156: 32'b01111011010100110101000010001000;
		10'd157: 32'b00110000000010001010000011101110;
		10'd158: 32'b11110101110010011100011000011100;
		10'd159: 32'b00110000110101000000100100101001;
		10'd160: 32'b00101110101111100101100001100000;
		10'd161: 32'b10011000100000010001101010011010;
		10'd162: 32'b00110100100100000000011000000000;
		10'd163: 32'b00011111000001100011000101000010;
		10'd164: 32'b01000011111101001000101111101010;
		10'd165: 32'b10101000100100000001111000000101;
		10'd166: 32'b01110001100000000010000001101100;
		10'd167: 32'b10010111110000010011100100000010;
		10'd168: 32'b01100100110000100010000101000110;
		10'd169: 32'b00011100010011000000011010000100;
		10'd170: 32'b10001000100010000010011000010100;
		10'd171: 32'b00000001000001010101011110011010;
		10'd172: 32'b00101100000110001000110010110100;
		10'd173: 32'b00000100001011111001010010000001;
		10'd174: 32'b00010001100011010000111001011100;
		10'd175: 32'b01110101000100000000101100100010;
		10'd176: 32'b11010000000010100010111001110000;
		10'd177: 32'b11010011010011000000101110100001;
		10'd178: 32'b00000100000000000000010111011001;
		10'd179: 32'b01010101000100000000000001011000;
		10'd180: 32'b11000110101001000101011010111000;
		10'd181: 32'b00101110001110000001100110000110;
		10'd182: 32'b10011011101000010001001010110000;
		10'd183: 32'b01110010000000001011000010100110;
		10'd184: 32'b00000110101101110100110001101101;
		10'd185: 32'b01100000101101000000111100011001;
		10'd186: 32'b01100000100001011000100110001110;
		10'd187: 32'b01010010001010011000001000100100;
		10'd188: 32'b00010000110101111101011000010101;
		10'd189: 32'b10010000000110101000011100100010;
		10'd190: 32'b01100100100101100000110110010010;
		10'd191: 32'b01001100010110101001001110011001;
		10'd192: 32'b01000001001100001100000010001101;
		10'd193: 32'b00000010011110010101111001000001;
		10'd194: 32'b00000100000001000011101010100010;
		10'd195: 32'b00000010101100010010111000000111;
		10'd196: 32'b01100100010000000000110000011101;
		10'd197: 32'b00101001011110001001000001010010;
		10'd198: 32'b00110101000010001000000101001100;
		10'd199: 32'b00100010010110010000000101000011;
		10'd200: 32'b00001000001110100100010010000000;
		10'd201: 32'b01100000100001001110000110011101;
		10'd202: 32'b00110101010101000110010001000101;
		10'd203: 32'b01000011110001010001000000010101;
		10'd204: 32'b01100010100110011010000101110000;
		10'd205: 32'b01110011110010010101100100010000;
		10'd206: 32'b01101100100001000100001011100001;
		10'd207: 32'b01101001010010101000000110101000;
		10'd208: 32'b01100011000001011010000011000010;
		10'd209: 32'b01001111000100100000110010101000;
		10'd210: 32'b00000110110110010010110011100000;
		10'd211: 32'b00011010110000111000001111000110;
		10'd212: 32'b00000011101100010000101010001010;
		10'd213: 32'b01001000110000100010000100101001;
		10'd214: 32'b00000001001001100000010001111001;
		10'd215: 32'b00000000111000011010010000100101;
		10'd216: 32'b10100101101000000111000010000110;
		10'd217: 32'b01100110011100101111001010001100;
		10'd218: 32'b00010000001011111010000001000010;
		10'd219: 32'b10000100111111101011010000011101;
		10'd220: 32'b00000100111001010010010111000000;
		10'd221: 32'b01111001011111001110100110011100;
		10'd222: 32'b10000000001001000010010010000110;
		10'd223: 32'b00111011101000110000010000000101;
		10'd224: 32'b10010100010000011000001000011010;
		10'd225: 32'b01001101000101111000100110100010;
		10'd226: 32'b10010001100111100101000110100100;
		10'd227: 32'b00000111000101111011001110000000;
		10'd228: 32'b10011110000010001001100100010110;
		10'd229: 32'b10101010000010010100100110001000;
		10'd230: 32'b11011000111000010100001110110000;
		10'd231: 32'b00100011101100101001010001000010;
		10'd232: 32'b00100001001100000111101000100010;
		10'd233: 32'b10000001100101010010011110101110;
		10'd234: 32'b01100100000010001111000010001011;
		10'd235: 32'b00010100000100100000100000101000;
		10'd236: 32'b00111100101100001000100001101010;
		10'd237: 32'b10001001110100010001111101011100;
		10'd238: 32'b10100000100110000100001011101000;
		10'd239: 32'b00001101101000100111100110111000;
		10'd240: 32'b00001000000000110100111100001010;
		10'd241: 32'b10111000110100000001010111110100;
		10'd242: 32'b10001101000101111010100110000000;
		10'd243: 32'b01001101100010000101101110000011;
		10'd244: 32'b00000000000101011110001110010001;
		10'd245: 32'b11000001101100010101100110100100;
		10'd246: 32'b00111100100000000011110010001010;
		10'd247: 32'b10000011100000100011100010011010;
		10'd248: 32'b01110100101010110000000110101011;
		10'd249: 32'b01010000000001101011000010011100;
		10'd250: 32'b10010011101101110000000001000001;
		10'd251: 32'b00010100000000110001001110000100;
		10'd252: 32'b01100010010000110000000011101011;
		10'd253: 32'b01000000000011010000000110011000;
		10'd254: 32'b01000011011000100001010111011000;
		10'd255: 32'b01000100010111001010010101000000;
		10'd256: 32'b11001000110000001111110110011101;
		10'd257: 32'b11000000010100101110010101010010;
		10'd258: 32'b11001001100000100011010000000000;
		10'd259: 32'b01001010011100001110101101000000;
		10'd260: 32'b10001011100000100101010111001101;
		10'd261: 32'b01010110010101110110110000111000;
		10'd262: 32'b00000001110000000011011110110100;
		10'd263: 32'b00111001101101000001111001101100;
		10'd264: 32'b01110101010101101100110010010000;
		10'd265: 32'b10001000110100100001100000011011;
		10'd266: 32'b01001001010000000000110011010001;
		10'd267: 32'b00110000000101100010011100010010;
		10'd268: 32'b10101101110101100101000010011011;
		10'd269: 32'b10000000010100100111100010110111;
		10'd270: 32'b00110000001101001000110001101111;
		10'd271: 32'b00100110110100010100100100001010;
		10'd272: 32'b00001101011011100110000100001100;
		10'd273: 32'b01100100100011000101010000100010;
		10'd274: 32'b01000101011100101001010001000000;
		10'd275: 32'b01110111110001001101110101110010;
		10'd276: 32'b11110101011010001001000100011000;
		10'd277: 32'b00100010110011101000101000000011;
		10'd278: 32'b01010101110001000101000000000000;
		10'd279: 32'b11011100001110100000111100010010;
		10'd280: 32'b01010101001010011001010111010001;
		10'd281: 32'b10110111101101000000000000000001;
		10'd282: 32'b11100101000100000010101110010000;
		10'd283: 32'b11001101001110110010011011110100;
		10'd284: 32'b11001110101010001000000010010000;
		10'd285: 32'b10001000101011011100100111111000;
		10'd286: 32'b11000010110010011000101010010000;
		10'd287: 32'b00100001010100001010110000100001;
		10'd288: 32'b10111000101100001111011010000101;
		10'd289: 32'b10001001110000001001010100000000;
		10'd290: 32'b01110001011100011010111001000011;
		10'd291: 32'b01011011110100110010000110010000;
		10'd292: 32'b10110101011100101010010000000011;
		10'd293: 32'b01011010010101101011110111000001;
		10'd294: 32'b10000101001100100010001101110100;
		10'd295: 32'b00101000011011000011110110101011;
		10'd296: 32'b00010100011010100101011110100110;
		10'd297: 32'b01010000110001100000011101010001;
		10'd298: 32'b11000010000011001001001010100100;
		10'd299: 32'b00010010000001000100110110000100;
		10'd300: 32'b11000010001010110010000000100000;
		10'd301: 32'b00000101101011001101100100000000;
		10'd302: 32'b11000011110011000100000110110000;
		10'd303: 32'b10101100110011100100110000100000;
		10'd304: 32'b10010000000010101001000100000100;
		10'd305: 32'b00000011110001011111100110000000;
		10'd306: 32'b00101100010000110100001000001101;
		10'd307: 32'b01101100100001100100001100010110;
		10'd308: 32'b00100001001001000000111000000100;
		10'd309: 32'b01010101010101110010101000001000;
		10'd310: 32'b01101100010001100000101000111111;
		10'd311: 32'b01100010001001001011000110100000;
		10'd312: 32'b01000001001000100100010010101110;
		10'd313: 32'b10001001001101110001100011000000;
		10'd314: 32'b10011000010000101011100000001010;
		10'd315: 32'b01110110010001000100000010000110;
		10'd316: 32'b01110000110101010001000010000001;
		10'd317: 32'b01100011101100011011000110000010;
		10'd318: 32'b10011010011010010000010000001000;
		10'd319: 32'b00000110111000100001010110010001;
		10'd320: 32'b11001001001000110111001100000000;
		10'd321: 32'b10000101011010111111001100111100;
		10'd322: 32'b00011110101110100000011100000000;
		10'd323: 32'b11110110111000010011100000000000;
		10'd324: 32'b00011010001000100110101100010100;
		10'd325: 32'b01000000111110010000000101110100;
		10'd326: 32'b10010111111110110111010000100000;
		10'd327: 32'b10100101101010101000001010110001;
		10'd328: 32'b00000000011011011010011100000111;
		10'd329: 32'b00101111001100000000000011111100;
		10'd330: 32'b00000001110010011100010101010101;
		10'd331: 32'b00100011101000011001101001001001;
		10'd332: 32'b11100100111111011010111101000010;
		10'd333: 32'b00111001100010000111010101001111;
		10'd334: 32'b10110101011001010001000100001001;
		10'd335: 32'b10110001010100010000111001001001;
		10'd336: 32'b00100100010001000000100100100100;
		10'd337: 32'b00011111010000000110010000001011;
		10'd338: 32'b11001000101000000000010010001111;
		10'd339: 32'b10110001010110010101101001001011;
		10'd340: 32'b00000001101110000110100100011011;
		10'd341: 32'b10111010010000000011010001101100;
		10'd342: 32'b11000101001000000010110100100011;
		10'd343: 32'b11011110110110001110100100000001;
		10'd344: 32'b10111011010101110100000010111000;
		10'd345: 32'b10001001010111110010110000000011;
		10'd346: 32'b10100001001000000100100110100001;
		10'd347: 32'b11001000110010011000101000010001;
		10'd348: 32'b00100000011110001100010110100000;
		10'd349: 32'b00000011110010110100010000001111;
		10'd350: 32'b00000001011010000100000000000101;
		10'd351: 32'b11100100001011001010001010001001;
		10'd352: 32'b00100111100101110111000010110000;
		10'd353: 32'b11001001111010010010000110001000;
		10'd354: 32'b00110000110000000010110011101100;
		10'd355: 32'b00101110010010010000101000101011;
		10'd356: 32'b00011001101000010000000011000001;
		10'd357: 32'b00001010010000110001001110101001;
		10'd358: 32'b10000110100001011010001000111101;
		10'd359: 32'b11101001000000101001011110101000;
		10'd360: 32'b10000010000110101110011010100000;
		10'd361: 32'b01000010000100001000010010000000;
		10'd362: 32'b00011110000001001111011000001000;
		10'd363: 32'b10011000001100001010010100100101;
		10'd364: 32'b00000111000110001000001000101010;
		10'd365: 32'b01001101111000110110000000101110;
		10'd366: 32'b01000110100111001110000001000100;
		10'd367: 32'b10101000101011101100001110110001;
		10'd368: 32'b01011110110100101000000011000000;
		10'd369: 32'b01111101001011010111000000000000;
		10'd370: 32'b00000011000101001001011100101111;
		10'd371: 32'b00100001001010110010101110100101;
		10'd372: 32'b11001100110100100001000001100100;
		10'd373: 32'b11110001010101000110110010100001;
		10'd374: 32'b10000110000000000001001111100110;
		10'd375: 32'b10000001100000100111011011110111;
		10'd376: 32'b00110101101100100100001011001111;
		10'd377: 32'b01011101101110000011000101110101;
		10'd378: 32'b00111001100010000001101011110100;
		10'd379: 32'b01001000110010000001000011110100;
		10'd380: 32'b00111001001010000101110001010011;
		10'd381: 32'b00111100001000110010010001010011;
		10'd382: 32'b00111100001100010011001011110110;
		10'd383: 32'b10010111000001100001010100100000;
		10'd384: 32'b00011111010101011110001001011100;
		10'd385: 32'b10100111010110101010100001111000;
		10'd386: 32'b01000100000010010111001000001010;
		10'd387: 32'b10011101001000001011011101110011;
		10'd388: 32'b10011111011000100000010001010000;
		10'd389: 32'b10100101100010000010010110111010;
		10'd390: 32'b11100010011010000101000000000010;
		10'd391: 32'b01101100000000001011100011001001;
		10'd392: 32'b01100010100100100100000100000010;
		10'd393: 32'b01000011010100001010010000101110;
		10'd394: 32'b11000000011100000101001011011010;
		10'd395: 32'b01111011100010101000110010001100;
		10'd396: 32'b10101100010011110101001101000110;
		10'd397: 32'b11100110110000000101001100000010;
		10'd398: 32'b00100011111110001100011000001010;
		10'd399: 32'b01010110011001110000010000100101;
		10'd400: 32'b10000100010000000110110100100110;
		10'd401: 32'b01000011010000100000100000111001;
		10'd402: 32'b00000010010100001000000010111101;
		10'd403: 32'b01000011000000100100011000111000;
		10'd404: 32'b10000000111000110011010010010111;
		10'd405: 32'b11110111010110110010011001111000;
		10'd406: 32'b00010101110010000110001001110110;
		10'd407: 32'b10001000100100110011000111100000;
		10'd408: 32'b00010110100110100101001011100101;
		10'd409: 32'b00101100100111110100110111000100;
		10'd410: 32'b00001000000100100000111010000000;
		10'd411: 32'b01111000000100100100111000010001;
		10'd412: 32'b10111110111110101011010011001101;
		10'd413: 32'b00011111000110010000000101000101;
		10'd414: 32'b10010100101000011000110110000001;
		10'd415: 32'b00110110001000000110001000000000;
		10'd416: 32'b10000010000111100000011011110001;
		10'd417: 32'b10011011010100100010000001000100;
		10'd418: 32'b11001001111011100011001110011001;
		10'd419: 32'b11101010000000010111110101010100;
		10'd420: 32'b01110000001011100101010010110111;
		10'd421: 32'b00001000000000100010010101000010;
		10'd422: 32'b10011100101011100001110000011110;
		10'd423: 32'b10011011011000100110000010010000;
		10'd424: 32'b10101000000001010000000100010110;
		10'd425: 32'b11110000000000010000100110110100;
		10'd426: 32'b01100100100011010011011110000010;
		10'd427: 32'b10000000101101010000000010000001;
		10'd428: 32'b00110000101011010000100100101000;
		10'd429: 32'b10111001101100011000000000000100;
		10'd430: 32'b11000100101111010001111100010111;
		10'd431: 32'b11110111001000010011000100101000;
		10'd432: 32'b10000010100000000111011011000110;
		10'd433: 32'b00100101001101000110000011000010;
		10'd434: 32'b11101110001000000100101100001100;
		10'd435: 32'b11010000100101000100001100000000;
		10'd436: 32'b00000010011000010111011100000001;
		10'd437: 32'b00110000010100000011101010101001;
		10'd438: 32'b11000010110000000111111000011000;
		10'd439: 32'b10000101111011011000110010001010;
		10'd440: 32'b10011001000101100001011000010011;
		10'd441: 32'b01001101000010001000101001100110;
		10'd442: 32'b00001100000000100011011100100100;
		10'd443: 32'b11010110001110110000110000010010;
		10'd444: 32'b00010000000110101101010000010101;
		10'd445: 32'b00010001101000001000000000100010;
		10'd446: 32'b01011000000110010011010111000110;
		10'd447: 32'b10000000001100010001101000100100;
		10'd448: 32'b00010000101010011110101101001111;
		10'd449: 32'b01111110001000010111100010000101;
		10'd450: 32'b00100010000110100110101000011000;
		10'd451: 32'b00100001100011011111111010110001;
		10'd452: 32'b10100001111000100101001011111010;
		10'd453: 32'b00010010011000000100101010000001;
		10'd454: 32'b11110000100010001011101000001010;
		10'd455: 32'b00001011001000000010100000110111;
		10'd456: 32'b00001000001100000100100100000001;
		10'd457: 32'b01000010111101001101000110111011;
		10'd458: 32'b11001000000000001100100010011000;
		10'd459: 32'b00101111100000011011101010010100;
		10'd460: 32'b10001010001111111000101100000001;
		10'd461: 32'b11000010001000000010110101010011;
		10'd462: 32'b00011000000000000011100000010000;
		10'd463: 32'b00100001000001000100011000001000;
		10'd464: 32'b00100100011110001100100000000000;
		10'd465: 32'b00000000001010001000000010011001;
		10'd466: 32'b10010011111011101100110011011010;
		10'd467: 32'b00100100010010101011010001011110;
		10'd468: 32'b00000101100000001000010000001000;
		10'd469: 32'b00000100011010000100110000001000;
		10'd470: 32'b11110101011011010000000111001011;
		10'd471: 32'b00101110000000100010011100100000;
		10'd472: 32'b01111101001010100110010000110000;
		10'd473: 32'b00100001010010000010100010011001;
		10'd474: 32'b00011001100001000110111000100001;
		10'd475: 32'b01000011000100111110001000100100;
		10'd476: 32'b01000110010001110101000001110000;
		10'd477: 32'b01101001010001001010101001110000;
		10'd478: 32'b00001011010000000110011000101100;
		10'd479: 32'b00110010000010000100001010000000;
		10'd480: 32'b01100010011000000010000101110000;
		10'd481: 32'b10101110001000001100101110000010;
		10'd482: 32'b01100100010000111010001011000011;
		10'd483: 32'b01010000011011000100110010110101;
		10'd484: 32'b10100000101011001100101000010110;
		10'd485: 32'b01101000100000101100101011011000;
		10'd486: 32'b00000000001101000000110100001100;
		10'd487: 32'b10110001001100001000011000101101;
		10'd488: 32'b00100010111000000000011101100010;
		10'd489: 32'b11100001001001110000001000001000;
		10'd490: 32'b00010000111011111001000001000011;
		10'd491: 32'b10101100110000011000011101101111;
		10'd492: 32'b00101010101000101000000000100110;
		10'd493: 32'b00000000011011001000100000011100;
		10'd494: 32'b10101000110000011001110010000011;
		10'd495: 32'b00000101001101010010010100010001;
		10'd496: 32'b10000010001000100100001000100110;
		10'd497: 32'b00110000001010010000011000010100;
		10'd498: 32'b00111000111100100001001000110101;
		10'd499: 32'b00010001010011000110101000010001;
		10'd500: 32'b10110100001000001111000001101100;
		10'd501: 32'b01000010110010111000010010001000;
		10'd502: 32'b00100111001010000010101000011100;
		10'd503: 32'b01001100100101001000100010111111;
		10'd504: 32'b00001111101001111010001111000110;
		10'd505: 32'b10000001101000110001100000000011;
		10'd506: 32'b10100011011110110001000110001011;
		10'd507: 32'b11001110000000110000110000010010;
		10'd508: 32'b00011100100010000000111100000001;
		10'd509: 32'b11100000010100011001000000000001;
		10'd510: 32'b10101010001101100110000100101101;
		10'd511: 32'b01100100011001100000011001001001;
		10'd512: 32'b01000101001000110000110011100010;
		10'd513: 32'b01001011000101010010001100101111;
		10'd514: 32'b11010001001101011001101010111000;
		10'd515: 32'b11100101001001010001010110001110;
		10'd516: 32'b01011000101101110010100110000110;
		10'd517: 32'b01101001100000000100001110000010;
		10'd518: 32'b11110111000101110010100000010001;
		10'd519: 32'b10111101101010000010100001000111;
		10'd520: 32'b10110001100001000001001000101100;
		10'd521: 32'b10101100001011000000000001111000;
		10'd522: 32'b11010101101100101100111000110011;
		10'd523: 32'b00001010110000011100101001100001;
		10'd524: 32'b01011110000111000011100000011110;
		10'd525: 32'b01011000001001111110100100010011;
		10'd526: 32'b11100000101100000100100100100000;
		10'd527: 32'b00100011000011000001000000010110;
		10'd528: 32'b11110011010000101001000111111010;
		10'd529: 32'b11010001000001010110101000011010;
		10'd530: 32'b10100000001101000001100100000010;
		10'd531: 32'b11000001100010000001001001100010;
		10'd532: 32'b01101101011001000101001111010010;
		10'd533: 32'b01011000001101110011010010111011;
		10'd534: 32'b10101001001111101000100111010110;
		10'd535: 32'b10000001100000101011111000100110;
		10'd536: 32'b00010001010001001111100010011110;
		10'd537: 32'b10000010011111101001000000100000;
		10'd538: 32'b00000110001011010010110010110001;
		10'd539: 32'b11100001000111001010010000100100;
		10'd540: 32'b00110010011000000010101010110100;
		10'd541: 32'b10010000011001001110011010010001;
		10'd542: 32'b00001000011000000111110011101111;
		10'd543: 32'b01110000101010001000001001000110;
		10'd544: 32'b00000010010100010110101101110100;
		10'd545: 32'b10100010000100011010010010110001;
		10'd546: 32'b00100101110100000001001001000100;
		10'd547: 32'b00010000010011000000100010000000;
		10'd548: 32'b00000100100101001010100001000100;
		10'd549: 32'b00010101000101000011110100010010;
		10'd550: 32'b00000011110001011001001001000101;
		10'd551: 32'b00101011001110010100110000001000;
		10'd552: 32'b10101011111000101101000110000110;
		10'd553: 32'b00000000111110110010100100111000;
		10'd554: 32'b11100000010110001010010110100000;
		10'd555: 32'b00011001001000010101110000110101;
		10'd556: 32'b00000111101110100110100111000101;
		10'd557: 32'b01000010110111001100111001111101;
		10'd558: 32'b11011001000100010100010001001100;
		10'd559: 32'b01111000110010000011100001010100;
		10'd560: 32'b01001010001100100100001001010010;
		10'd561: 32'b01010011111100001000000111101001;
		10'd562: 32'b00101000100101111000101011001001;
		10'd563: 32'b01101000101011111010100111001000;
		10'd564: 32'b00101000101100100000000001000000;
		10'd565: 32'b00001111010000010001000001001101;
		10'd566: 32'b00101000001000110000100001110110;
		10'd567: 32'b00100101010000000000010000010100;
		10'd568: 32'b01111010100001110001100111000000;
		10'd569: 32'b10111111110010011101100100000100;
		10'd570: 32'b01101001011000010001110101000110;
		10'd571: 32'b10000101111101000000000010100100;
		10'd572: 32'b00100011000010000001010011110010;
		10'd573: 32'b00111101100001101110010111001000;
		10'd574: 32'b01001010100000010101111010000100;
	endcase;
	return out;
endfunction
function Bit#(32) get_output_page3(UInt#(10) counter);
	Bit#(32) out = case(counter)
		10'd0: 32'b01000100100010000100010010001000;
		10'd1: 32'b00010000000101000000000000110100;
		10'd2: 32'b00000100001000000000000001100010;
		10'd3: 32'b00000011000000100000001101010010;
		10'd4: 32'b00000100001000000100000001100000;
		10'd5: 32'b10000000000100010000000000010000;
		10'd6: 32'b01000000000010100100000100010010;
		10'd7: 32'b00000000000000110001000101000110;
		10'd8: 32'b00000100000000000010000101000010;
		10'd9: 32'b00000101001001010000010000010101;
		10'd10: 32'b00010001000000010000000000000110;
		10'd11: 32'b00010001000100000000000000010010;
		10'd12: 32'b00000000010100000000000101100000;
		10'd13: 32'b00000000101000100000000000110100;
		10'd14: 32'b00000100001101000000010000100000;
		10'd15: 32'b01000000000000000111000100000000;
		10'd16: 32'b00011000010000110001100000000011;
		10'd17: 32'b11100000000001100110000000000110;
		10'd18: 32'b00010000000000010000001010000001;
		10'd19: 32'b00000000000000010101000010000111;
		10'd20: 32'b00000000000011100000000000010011;
		10'd21: 32'b00000100101000010000000000001100;
		10'd22: 32'b00010000000100010000000100010010;
		10'd23: 32'b01100000000000000000000000101000;
		10'd24: 32'b01000000000000010100000100000010;
		10'd25: 32'b00100000001000010010000000100000;
		10'd26: 32'b00110000000100000010000000010000;
		10'd27: 32'b00000000110100100000000111000010;
		10'd28: 32'b00000011000000100001000100000110;
		10'd29: 32'b00010100000100110001000000000000;
		10'd30: 32'b00010001001000100001000100100110;
		10'd31: 32'b10000000000100001000010000001000;
		10'd32: 32'b10010000110000001001000000010000;
		10'd33: 32'b01000100010000000000001001010000;
		10'd34: 32'b00110000000000001100000000001010;
		10'd35: 32'b00000001000100100000000100010101;
		10'd36: 32'b01000000010100000000000001010010;
		10'd37: 32'b00000000011000000001000001110000;
		10'd38: 32'b00010010000000100001001000000100;
		10'd39: 32'b00100000000010000000010000000010;
		10'd40: 32'b00011000100000010000100000000010;
		10'd41: 32'b00000010000000111100000000000110;
		10'd42: 32'b01000000000100100000000000100110;
		10'd43: 32'b00000000000000010110001000100001;
		10'd44: 32'b00100000000000010010000100010001;
		10'd45: 32'b00000001000100000000001100000010;
		10'd46: 32'b00001000010000010010000001000000;
		10'd47: 32'b11000100000010000000000000100000;
		10'd48: 32'b00000000100100000000000101010000;
		10'd49: 32'b10100000000001001011000000000000;
		10'd50: 32'b01010000000000110000010100000110;
		10'd51: 32'b00000001010000010100000100000001;
		10'd52: 32'b10000100000000101000010100000001;
		10'd53: 32'b00000101000001000000011000000110;
		10'd54: 32'b01010000000101000100000000000110;
		10'd55: 32'b00011000000000000001100000001001;
		10'd56: 32'b00000000100100000000000011010101;
		10'd57: 32'b00100001000000110000000100000001;
		10'd58: 32'b00010000010000010000010001000010;
		10'd59: 32'b10000000000001100000000000000110;
		10'd60: 32'b00100000000000100001000100000110;
		10'd61: 32'b00000000100001000010000010000000;
		10'd62: 32'b01000010000000010000001000010001;
		10'd63: 32'b11110011000110111010110110001001;
		10'd64: 32'b11101111110111101100010100101000;
		10'd65: 32'b11100000110110101010010101101111;
		10'd66: 32'b11111101110001001001000101001101;
		10'd67: 32'b11000011011110110111010101000000;
		10'd68: 32'b01110011111111101100100011010100;
		10'd69: 32'b01010101100010100110100101110000;
		10'd70: 32'b10100111100000111011011101101011;
		10'd71: 32'b00111110010010010101001000001001;
		10'd72: 32'b11000101100110011000110100101011;
		10'd73: 32'b11000101001001010110011101001100;
		10'd74: 32'b11110011000101110001001000001010;
		10'd75: 32'b10000101001000110010011110000000;
		10'd76: 32'b10111100010010010111001110001001;
		10'd77: 32'b10000001000011000001001101011000;
		10'd78: 32'b11110101011101101111001110101111;
		10'd79: 32'b11101010011000111110111101110001;
		10'd80: 32'b01010110000101011100011001101011;
		10'd81: 32'b00001110111010101111110011000110;
		10'd82: 32'b01010001011100000011011000100100;
		10'd83: 32'b11011010111101001101001000110010;
		10'd84: 32'b01100110000010110111110101001001;
		10'd85: 32'b10011010011010100001110001111101;
		10'd86: 32'b11000000001110100011011001100110;
		10'd87: 32'b00101100001011011010100111010101;
		10'd88: 32'b10011101101011111110100111010001;
		10'd89: 32'b01000111010111010011001010100101;
		10'd90: 32'b11110001001111100011001110000110;
		10'd91: 32'b00100101000010000010011001010011;
		10'd92: 32'b01000111111101100000101101101011;
		10'd93: 32'b00110101010101001100111100110011;
		10'd94: 32'b01000010101001000001111101010111;
		10'd95: 32'b01101101010111010010010111001011;
		10'd96: 32'b00011000000101010101000000001001;
		10'd97: 32'b10001111010101011000110010001111;
		10'd98: 32'b10110100101011110101011100000111;
		10'd99: 32'b11000100010010010110110000000101;
		10'd100: 32'b01101110111001010110001000001000;
		10'd101: 32'b11000001010001110000011100001011;
		10'd102: 32'b00111101000000011001000101000001;
		10'd103: 32'b10101111100000100011001010001101;
		10'd104: 32'b11010111110101111110000100111100;
		10'd105: 32'b10011111011101101000010110110010;
		10'd106: 32'b00000011111110100110100010010011;
		10'd107: 32'b00101111110101111000001110001100;
		10'd108: 32'b11011111111101011011111100011000;
		10'd109: 32'b00001011111010101101000101010101;
		10'd110: 32'b01011010100010101100011001101001;
		10'd111: 32'b00111100111011111111011011111010;
		10'd112: 32'b11110101000101100110001101110111;
		10'd113: 32'b00000100010100000111101000110011;
		10'd114: 32'b11110011000111101100111001101011;
		10'd115: 32'b00110110000011111101001011100111;
		10'd116: 32'b11100010111001001010010000111001;
		10'd117: 32'b10011010000111100111001011010110;
		10'd118: 32'b11011001001111101000101011110011;
		10'd119: 32'b00111000010100100001100001010110;
		10'd120: 32'b10010100100000011011010011110010;
		10'd121: 32'b01110110000100100001100000011111;
		10'd122: 32'b10100101010100100001010011101101;
		10'd123: 32'b00111110000000000011101011010010;
		10'd124: 32'b00011100010001011000100100110111;
		10'd125: 32'b00110111011110000100110100010110;
		10'd126: 32'b11111011100100010100110110111011;
		10'd127: 32'b01111011001010001111101110010001;
		10'd128: 32'b01111010110100111100010000000010;
		10'd129: 32'b00100010011111000111001010011101;
		10'd130: 32'b01100111101110101010000111110111;
		10'd131: 32'b01001111001010000100000101111011;
		10'd132: 32'b10011001101101001110100010000010;
		10'd133: 32'b00100100101011000001100011011100;
		10'd134: 32'b11111011011111101111100101011111;
		10'd135: 32'b10111101011000011000100111101000;
		10'd136: 32'b11111101000100111110100000100010;
		10'd137: 32'b11000101110001111000100000001101;
		10'd138: 32'b11111111110111101001100110000101;
		10'd139: 32'b10001100100000000011110000101010;
		10'd140: 32'b00111010100110001000101101111000;
		10'd141: 32'b00111111010000111111111110001101;
		10'd142: 32'b11101111110011100001101110001000;
		10'd143: 32'b00111100001100010100010000010010;
		10'd144: 32'b11000010111011001000100010111111;
		10'd145: 32'b00101100100100100111111001001001;
		10'd146: 32'b11111101111010111100100010101001;
		10'd147: 32'b00100100001011001101111100010001;
		10'd148: 32'b00111000010101010110100011100111;
		10'd149: 32'b10100010010000011111011101010000;
		10'd150: 32'b10111010111010000110100011101000;
		10'd151: 32'b10000101100001000110000110001000;
		10'd152: 32'b11001111111111011010010110000000;
		10'd153: 32'b00101000100011111010000000001010;
		10'd154: 32'b11110001110001011010100110111000;
		10'd155: 32'b00101011101101000110010110011011;
		10'd156: 32'b01111011010100110101000010001000;
		10'd157: 32'b01110001000010001110000011101110;
		10'd158: 32'b11111101110010011100011010011100;
		10'd159: 32'b00110000110101110001100100111001;
		10'd160: 32'b01111110101111100101101001110000;
		10'd161: 32'b10011000100101010001101010011010;
		10'd162: 32'b11110111100101000000011100110100;
		10'd163: 32'b00011111100001100011001101000010;
		10'd164: 32'b11000111111111001000101111101010;
		10'd165: 32'b11101000100100000001111000010101;
		10'd166: 32'b01110001100010000110001001101100;
		10'd167: 32'b10010111110001110011100100011110;
		10'd168: 32'b01100100110010110010010111000111;
		10'd169: 32'b00011100011011000000011010000100;
		10'd170: 32'b10001001100011000010011100010100;
		10'd171: 32'b01001001000001010101111110111110;
		10'd172: 32'b00101100100110001000110010110100;
		10'd173: 32'b00001100001011111001010010000111;
		10'd174: 32'b01010001100111010011111001011100;
		10'd175: 32'b01110101000100010000101101100011;
		10'd176: 32'b11010000000010100011111001111000;
		10'd177: 32'b11010111011111000000111110111101;
		10'd178: 32'b00000110000000000000011111011001;
		10'd179: 32'b01010111000101000000001011011001;
		10'd180: 32'b11000110111001000101011010111010;
		10'd181: 32'b00101110011111000001100110000110;
		10'd182: 32'b10011011101000010011001010110000;
		10'd183: 32'b01110110000000001011000010100110;
		10'd184: 32'b10001110101101110100111001101101;
		10'd185: 32'b11110001101101010000111100111001;
		10'd186: 32'b01110000100001011000100110001110;
		10'd187: 32'b01110010001010011000001001100100;
		10'd188: 32'b00010000110111111101111110110101;
		10'd189: 32'b10010000001110101000011110100010;
		10'd190: 32'b01110110101101100000110110110110;
		10'd191: 32'b01001100010110101001001110011101;
		10'd192: 32'b01000001001100001101000010001101;
		10'd193: 32'b00000011011110010101111001101011;
		10'd194: 32'b01011100000001000011101110100110;
		10'd195: 32'b00000010101100110110111000001111;
		10'd196: 32'b01100100110100000000110000011101;
		10'd197: 32'b10111001011110101001000001010011;
		10'd198: 32'b00111101000010101000000101101100;
		10'd199: 32'b00100010010111010101010101000011;
		10'd200: 32'b00001000001111100100011011000000;
		10'd201: 32'b01100000110001001110010110011101;
		10'd202: 32'b01110101010101000110010001000101;
		10'd203: 32'b01010011110001010101010001010101;
		10'd204: 32'b11101110100110011010000101110001;
		10'd205: 32'b01110011110010010111110100011001;
		10'd206: 32'b01101101100001000110001011100111;
		10'd207: 32'b01111001010010101000010110101000;
		10'd208: 32'b01100011001001011010001011000110;
		10'd209: 32'b01001111000101100000110110101100;
		10'd210: 32'b00010110110110010010110011100000;
		10'd211: 32'b11011010110000111000001111000110;
		10'd212: 32'b00000111101100010001101110011011;
		10'd213: 32'b01001010110100100010000110101001;
		10'd214: 32'b00000001001001100011010001111001;
		10'd215: 32'b10000000111001011110010000111101;
		10'd216: 32'b10100101101000000111000010000110;
		10'd217: 32'b01100111011100101111001110001101;
		10'd218: 32'b00110100001011111010001001000010;
		10'd219: 32'b11010100111111101011011000011101;
		10'd220: 32'b00000101111001010010010111000000;
		10'd221: 32'b01111001011111001111110110111100;
		10'd222: 32'b10000100111001011010010010000110;
		10'd223: 32'b10111011101000110000011100100101;
		10'd224: 32'b10010100010000111000001100111110;
		10'd225: 32'b01011101011111111000100110100010;
		10'd226: 32'b10010001110111100101000110101100;
		10'd227: 32'b00000111000101111011101110000000;
		10'd228: 32'b10011110010010011001100100010110;
		10'd229: 32'b10101011001010010101100110101010;
		10'd230: 32'b11011010111000011101001110110001;
		10'd231: 32'b10100011101110111001110101000010;
		10'd232: 32'b10100001101100000111101000101010;
		10'd233: 32'b10000101110111011111111110101110;
		10'd234: 32'b01100100100011001111000111001111;
		10'd235: 32'b00110101001100100000110000101010;
		10'd236: 32'b10111100101100101001101001101010;
		10'd237: 32'b10001001110100010001111101011100;
		10'd238: 32'b10100000100110000100001111101000;
		10'd239: 32'b00001101111000100111100110111000;
		10'd240: 32'b00001000001000110100111110001010;
		10'd241: 32'b10111001110100000001010111110100;
		10'd242: 32'b10001111101101111010101111000000;
		10'd243: 32'b11001101100010000111101110101011;
		10'd244: 32'b00100010000101111110101111010001;
		10'd245: 32'b11000011101100011111100110100100;
		10'd246: 32'b00111101100000000011110010001010;
		10'd247: 32'b10001011100000110011101010111010;
		10'd248: 32'b11110101101010110000000110101011;
		10'd249: 32'b01010000000011101011011110011101;
		10'd250: 32'b10010011101101111000000011100001;
		10'd251: 32'b10010100010001110001101110001101;
		10'd252: 32'b11111011010100111000000011101011;
		10'd253: 32'b01100101000011010000100111011000;
		10'd254: 32'b01000011111000110001010111011001;
		10'd255: 32'b01000100010111001110010101001010;
		10'd256: 32'b11001100110000001111111111011101;
		10'd257: 32'b11000010010101101110010101010010;
		10'd258: 32'b11001001110000100011010010110010;
		10'd259: 32'b11001011011100011111111101000000;
		10'd260: 32'b10001011100000110101010111011101;
		10'd261: 32'b01010110010101110110110101111110;
		10'd262: 32'b01000101110000100111011110110100;
		10'd263: 32'b00111001101101100001111001101110;
		10'd264: 32'b01110101010101101100110010010011;
		10'd265: 32'b10101000111100100001101100011011;
		10'd266: 32'b01001001011000110110110011010001;
		10'd267: 32'b00111000000101100010011100010010;
		10'd268: 32'b10111101110101110101000010011011;
		10'd269: 32'b10000000010101100111100010110111;
		10'd270: 32'b00111000101101001000110001101111;
		10'd271: 32'b00100111110100110100100100011011;
		10'd272: 32'b00001101111111100110001100101100;
		10'd273: 32'b01100100101011000101010000100010;
		10'd274: 32'b01010111011100101001010011000000;
		10'd275: 32'b01110111110001001101110101110010;
		10'd276: 32'b11110101111010001001100100011000;
		10'd277: 32'b00100011110011101000101001001111;
		10'd278: 32'b01111101111101100111000000000000;
		10'd279: 32'b11011100011110110000111100010010;
		10'd280: 32'b11010101001011011001010111011011;
		10'd281: 32'b10110111101101010100101110010001;
		10'd282: 32'b11100101010100010011111110010000;
		10'd283: 32'b11001101001110110010011011110100;
		10'd284: 32'b11001110101010011000011010010001;
		10'd285: 32'b10001100101011011110100111111000;
		10'd286: 32'b11000111110010011000101010011000;
		10'd287: 32'b01100001011100101010110010111101;
		10'd288: 32'b10111010101100011111011010000101;
		10'd289: 32'b11011101111100001011010100010000;
		10'd290: 32'b11110001111100111010111001000011;
		10'd291: 32'b01111111110100110010000111110000;
		10'd292: 32'b10110101111100111011011000000011;
		10'd293: 32'b11111010010101101011110111000111;
		10'd294: 32'b11100101011110100010001101111101;
		10'd295: 32'b00111000011011000011110110101011;
		10'd296: 32'b10110100011110100111011110111110;
		10'd297: 32'b01010010110001101000011101010011;
		10'd298: 32'b11000010000011001001011010110100;
		10'd299: 32'b00010010100011000100110110000110;
		10'd300: 32'b11010010101010110010000000101000;
		10'd301: 32'b10000101111011001111100100000000;
		10'd302: 32'b11001111110011000101010110110000;
		10'd303: 32'b10101100111011110110111000110000;
		10'd304: 32'b10010001000010111001001111100110;
		10'd305: 32'b00011011111101011111100110000101;
		10'd306: 32'b00101101010000110110001001001111;
		10'd307: 32'b01101100110011100100001100010110;
		10'd308: 32'b10101101111001100000111100000100;
		10'd309: 32'b01010101010111111010101000001000;
		10'd310: 32'b01101100110001110010101000111111;
		10'd311: 32'b01100010001001001011010110100000;
		10'd312: 32'b01000001001000110110110010101111;
		10'd313: 32'b11001101001101110001110011010110;
		10'd314: 32'b10011000010000101011100010001010;
		10'd315: 32'b11110110010001011100110010000110;
		10'd316: 32'b01110000111101011001010010000011;
		10'd317: 32'b11100011101101111011000111000010;
		10'd318: 32'b10111010011010010000010001001000;
		10'd319: 32'b00000111111000100101010111010001;
		10'd320: 32'b11001011101001110111001100000000;
		10'd321: 32'b10011111011010111111001100111110;
		10'd322: 32'b00011111111110100100011100100001;
		10'd323: 32'b11110110111001010011100000000001;
		10'd324: 32'b00011111001100111110111101110100;
		10'd325: 32'b11001000111110010100000101110111;
		10'd326: 32'b11010111111110110111010000100001;
		10'd327: 32'b10101111111010111001111010110011;
		10'd328: 32'b10000101011011111010011100001111;
		10'd329: 32'b10101111001110100010000011111110;
		10'd330: 32'b00001001110010011100011111011101;
		10'd331: 32'b00100011101000011001111001001001;
		10'd332: 32'b11100100111111111010111101100011;
		10'd333: 32'b00111001101111000111010101001111;
		10'd334: 32'b11110101011101011001010111001001;
		10'd335: 32'b10111011010100011001111001011001;
		10'd336: 32'b00100100010001000000101100110100;
		10'd337: 32'b10011111010000000110110000001011;
		10'd338: 32'b11001000101000000000010110101111;
		10'd339: 32'b11110011010110010101101001001011;
		10'd340: 32'b10001001111110000111111101011011;
		10'd341: 32'b10111010010010000011011101101110;
		10'd342: 32'b11001101101000010010110100101011;
		10'd343: 32'b11011110110110001110101111101011;
		10'd344: 32'b10111011010101110100000010111100;
		10'd345: 32'b10001001110111110110111010100011;
		10'd346: 32'b10100001011000000100100111100101;
		10'd347: 32'b11001101110011111000111100011001;
		10'd348: 32'b10100000111111001100010110110000;
		10'd349: 32'b11000111110110110100010000001111;
		10'd350: 32'b10001001011010000100001000000101;
		10'd351: 32'b11101100001111001010001010101001;
		10'd352: 32'b00101111101101110111000011110000;
		10'd353: 32'b11011001111010010010010110101001;
		10'd354: 32'b01110000110000000010111011101100;
		10'd355: 32'b00101110110011010010101100101011;
		10'd356: 32'b00011001101001010000000011000001;
		10'd357: 32'b00001010010100110001001110101011;
		10'd358: 32'b10000110100001111010111000111101;
		10'd359: 32'b11101001000010101001011110101000;
		10'd360: 32'b11000010000110101110011010100000;
		10'd361: 32'b01000010000110011000010110010100;
		10'd362: 32'b00111111100001001111011000101001;
		10'd363: 32'b11011001001100001010011100111101;
		10'd364: 32'b00000111000110101001001100101010;
		10'd365: 32'b01001101111000111110000010101110;
		10'd366: 32'b11000111100111001110010001100100;
		10'd367: 32'b10101000101011101110001110111001;
		10'd368: 32'b01011110110100111101000011000000;
		10'd369: 32'b01111101101011010111001000000000;
		10'd370: 32'b00000011000101001001011100101111;
		10'd371: 32'b10100001101010111010101110101101;
		10'd372: 32'b11001100110101100001000101100100;
		10'd373: 32'b11111001010101000110110010100001;
		10'd374: 32'b11000110001000000001101111101111;
		10'd375: 32'b10000001100000100111011011111111;
		10'd376: 32'b00110101101100100101011011011111;
		10'd377: 32'b01011101101110100011100101111101;
		10'd378: 32'b00111001100010001011111011111100;
		10'd379: 32'b01011000111010000001000011110110;
		10'd380: 32'b00111001101010100101110101011011;
		10'd381: 32'b00111101001101110010010011010111;
		10'd382: 32'b00111101101101010011001011110110;
		10'd383: 32'b10011111010011100001010100110000;
		10'd384: 32'b11011111010101011111001001011110;
		10'd385: 32'b10100111010110101011110111111000;
		10'd386: 32'b11000110001010110111101000001010;
		10'd387: 32'b10011101001000001011011111110011;
		10'd388: 32'b10011111011000101000110101010001;
		10'd389: 32'b10100101100010011010010110111010;
		10'd390: 32'b11110011011010010101110000000111;
		10'd391: 32'b01101100010100001011100011011101;
		10'd392: 32'b01101110101100100100011100000010;
		10'd393: 32'b01100011110100001110010001101110;
		10'd394: 32'b11101001111100000101001011011010;
		10'd395: 32'b01111011100010101000110010001100;
		10'd396: 32'b10101100010111110101011111010110;
		10'd397: 32'b11101110111000001111011100001010;
		10'd398: 32'b00100011111110101100011010011010;
		10'd399: 32'b01010111111001110001010000100101;
		10'd400: 32'b10100100010000000111111110110110;
		10'd401: 32'b11010011010001100000110000111001;
		10'd402: 32'b01100010110100001000100011111101;
		10'd403: 32'b01000011000000100100011000111101;
		10'd404: 32'b10000110111000110011010011010111;
		10'd405: 32'b11110111010110110010111001111100;
		10'd406: 32'b10010101111010001110011001111111;
		10'd407: 32'b10001000100110110011001111110100;
		10'd408: 32'b00010110101110111111001111100101;
		10'd409: 32'b00101110100111110100110111000100;
		10'd410: 32'b01001011111100110000111010010010;
		10'd411: 32'b01111000100100101100111101010101;
		10'd412: 32'b10111110111110101011010011001101;
		10'd413: 32'b00011111000110111000000111100101;
		10'd414: 32'b10010100111100111001111110000001;
		10'd415: 32'b00111110001100000111001101001000;
		10'd416: 32'b10100010001111100001011011111001;
		10'd417: 32'b10011011011100100010001011000100;
		10'd418: 32'b11001001111111100011001111011001;
		10'd419: 32'b11101010100000010111110101010100;
		10'd420: 32'b01110000001111100101010010110111;
		10'd421: 32'b10111011101100100010011101000010;
		10'd422: 32'b10111100101011100101110001011110;
		10'd423: 32'b10111011011000100110000011010100;
		10'd424: 32'b10111001100001110000010100010110;
		10'd425: 32'b11111000010010010000100110110110;
		10'd426: 32'b01100101100011010011011110001010;
		10'd427: 32'b10011000101101110000010011000001;
		10'd428: 32'b00111001101011010000100100111000;
		10'd429: 32'b10111001101100011000010100000110;
		10'd430: 32'b11000100101111011001111100011111;
		10'd431: 32'b11110111001000010111001100101001;
		10'd432: 32'b10100110100000000111011011000110;
		10'd433: 32'b00100101001101000110000111010010;
		10'd434: 32'b11101111011100010100111100101101;
		10'd435: 32'b11110000100101000110001100000100;
		10'd436: 32'b00110010011001011111011100000011;
		10'd437: 32'b00110000010100001111101010101001;
		10'd438: 32'b11001010110000100111111001111000;
		10'd439: 32'b11000101111011011100110010001010;
		10'd440: 32'b10011001001101100001011000010111;
		10'd441: 32'b01001101001011101001101001100110;
		10'd442: 32'b10011100000010100011011100110100;
		10'd443: 32'b11011110001110111000110010010010;
		10'd444: 32'b00010000000110101101010000010111;
		10'd445: 32'b00011101101010101001100010100010;
		10'd446: 32'b01011100000110010011010111000110;
		10'd447: 32'b10000000011100010001101010100101;
		10'd448: 32'b10011110101010011111101101001111;
		10'd449: 32'b01111110101000010111111010001101;
		10'd450: 32'b00110010000110101110101010011010;
		10'd451: 32'b10111001110011111111111111110001;
		10'd452: 32'b10101011111000100111001111111111;
		10'd453: 32'b00010010011000010111101010000111;
		10'd454: 32'b11110001111010001111111000001010;
		10'd455: 32'b00001011101000001010100001110111;
		10'd456: 32'b00001000011100000110100100010001;
		10'd457: 32'b01000011111101001101000110111011;
		10'd458: 32'b11001010110010001100100010011000;
		10'd459: 32'b00101111101000011011101110110100;
		10'd460: 32'b10001010001111111000101100000001;
		10'd461: 32'b11001010001000000010110101110111;
		10'd462: 32'b00011011000000001011100000010000;
		10'd463: 32'b11100001000011000110011100001010;
		10'd464: 32'b00110100011110001100100000000000;
		10'd465: 32'b00110000101010001000000010111001;
		10'd466: 32'b10010011111011101100110011011011;
		10'd467: 32'b00100100010010101011011001111110;
		10'd468: 32'b10000111100010001110010000001000;
		10'd469: 32'b00100100111110000100110000001010;
		10'd470: 32'b11110101011011010000100111001011;
		10'd471: 32'b00111110000000100010111100110000;
		10'd472: 32'b01111101101110100110110000110001;
		10'd473: 32'b00100011010010000010100010111001;
		10'd474: 32'b00011001100101000110111000100001;
		10'd475: 32'b01010011000100111110001000100100;
		10'd476: 32'b01001110010001110111010001110100;
		10'd477: 32'b01111001010001001010101011110000;
		10'd478: 32'b00001011010001000110011000111101;
		10'd479: 32'b10110010000010001110011010000000;
		10'd480: 32'b01100010011101001010100101110000;
		10'd481: 32'b11101110001000001100101111000110;
		10'd482: 32'b01100100010100111010001011000011;
		10'd483: 32'b01111010011011000110111010111101;
		10'd484: 32'b10100000111111001101101001110110;
		10'd485: 32'b11101000100001101100101011011000;
		10'd486: 32'b00000010011101001010110100001100;
		10'd487: 32'b10110101001110011000111000101101;
		10'd488: 32'b00100010111000001000011101100010;
		10'd489: 32'b11110001001011111010001000001110;
		10'd490: 32'b00010000111011111001110001000011;
		10'd491: 32'b10101100111000111000011101101111;
		10'd492: 32'b00101110101001101000100000110110;
		10'd493: 32'b00000010111111001000101100111101;
		10'd494: 32'b10101100110000011001110010000011;
		10'd495: 32'b00010101101101010010010101111001;
		10'd496: 32'b11110010011100100101001000101110;
		10'd497: 32'b00110010001010110000011000011100;
		10'd498: 32'b00111010111110101101001000111101;
		10'd499: 32'b00010001010011010111101100010001;
		10'd500: 32'b10110100001001001111000001101100;
		10'd501: 32'b01000010110010111000010010001000;
		10'd502: 32'b10111111001010100110101010111100;
		10'd503: 32'b01001101100101011000111010111111;
		10'd504: 32'b00001111101001111010011111111111;
		10'd505: 32'b11000011101000110101100000010011;
		10'd506: 32'b10100011011110110101000110101011;
		10'd507: 32'b11001110000000110100110000010011;
		10'd508: 32'b00111100110110100000111100000001;
		10'd509: 32'b11100010010100011001010000010001;
		10'd510: 32'b10101110001101110110000100101101;
		10'd511: 32'b01100100011101100010011001111001;
		10'd512: 32'b01000101001000110000110011100010;
		10'd513: 32'b01111011010101010010001110101111;
		10'd514: 32'b11010011101101111101101110111000;
		10'd515: 32'b11101101001001010011110110101110;
		10'd516: 32'b01011000101101110010100110010111;
		10'd517: 32'b01101001100100000100111110000010;
		10'd518: 32'b11110111001101110011100000010001;
		10'd519: 32'b10111101101010001010100001001111;
		10'd520: 32'b10111001100001000001101000101100;
		10'd521: 32'b10101100001011100000001011111000;
		10'd522: 32'b11111101101100101100111100111111;
		10'd523: 32'b00011110110010011100101001100001;
		10'd524: 32'b01011110010111000011110010011110;
		10'd525: 32'b01011000001001111110111100011011;
		10'd526: 32'b11110101101111000100100100100100;
		10'd527: 32'b00110011000011000001010000010110;
		10'd528: 32'b11110011011000101001100111111010;
		10'd529: 32'b11010001000001010111101001011110;
		10'd530: 32'b10100011001101000001100100000010;
		10'd531: 32'b11100001100010000001001001110010;
		10'd532: 32'b01111101011001100101001111010010;
		10'd533: 32'b01011001001101110011010011111111;
		10'd534: 32'b11101001001111101001100111010110;
		10'd535: 32'b11001001110000101111111000100110;
		10'd536: 32'b01110101011001001111100010011110;
		10'd537: 32'b10001110011111101011100100100000;
		10'd538: 32'b00100110101011011010110010110101;
		10'd539: 32'b11100001100111001011011100100111;
		10'd540: 32'b10110110011001000110101011110100;
		10'd541: 32'b10110010011001101110011010010001;
		10'd542: 32'b10001000011000001111111011101111;
		10'd543: 32'b01110000111010001000001101000110;
		10'd544: 32'b00001011110100010110101101111101;
		10'd545: 32'b11100010100100011010010010110011;
		10'd546: 32'b00100101110101000001101001010100;
		10'd547: 32'b00110000011011000000100010000000;
		10'd548: 32'b00010100110101001010100001000100;
		10'd549: 32'b00010101000101000011110110010011;
		10'd550: 32'b00100011110001111001001001001101;
		10'd551: 32'b01101011011111010100110000111000;
		10'd552: 32'b10101011111100111111011110000111;
		10'd553: 32'b00000001111110111010100100111100;
		10'd554: 32'b11100000010110001010110110100001;
		10'd555: 32'b11011001001100110101110000110101;
		10'd556: 32'b00000111101111101110100111000101;
		10'd557: 32'b01100011110111001100111001111101;
		10'd558: 32'b11011011001100110100010011001110;
		10'd559: 32'b11111000110110010111100001010100;
		10'd560: 32'b11001010011101100100001011010010;
		10'd561: 32'b01010011111100011000000111101011;
		10'd562: 32'b00101000100101111101101011101001;
		10'd563: 32'b01111001111111111011100111001101;
		10'd564: 32'b00101000101100100100000011000000;
		10'd565: 32'b00001111010000010001000001001101;
		10'd566: 32'b00101100001010110000100011110110;
		10'd567: 32'b00100111011011000000010000110100;
		10'd568: 32'b01111011100001110001111111100001;
		10'd569: 32'b10111111110010011101110100010100;
		10'd570: 32'b01101001011000010001111111010110;
		10'd571: 32'b10110101111111100000000010100100;
		10'd572: 32'b00111011010010001001010111110010;
		10'd573: 32'b00111101110011101110010111001100;
		10'd574: 32'b01111010110000010101111011010100;
	endcase;
	return out;
endfunction
function Bit#(32) get_output_page4(UInt#(10) counter);
	Bit#(32) out = case(counter)
		10'd0: 32'b01000100100011000100010010001000;
		10'd1: 32'b00110000000101000001000000110100;
		10'd2: 32'b00001100001000000000000001100010;
		10'd3: 32'b00010011000000100000001101010010;
		10'd4: 32'b00000101001001000100000001100000;
		10'd5: 32'b10000000010100010000000000010000;
		10'd6: 32'b01010000000010100101000100011010;
		10'd7: 32'b00000010010000110001000101000110;
		10'd8: 32'b10000100100000000010000101000010;
		10'd9: 32'b01000101001001110000010000010101;
		10'd10: 32'b00010001000000010000000100000110;
		10'd11: 32'b00010001000100000000000000011010;
		10'd12: 32'b00000000010110000000000101100000;
		10'd13: 32'b00000000101000100000000000110101;
		10'd14: 32'b00000100001101100000010000100000;
		10'd15: 32'b01000000010000000111000101000000;
		10'd16: 32'b00011000010001110001110000000011;
		10'd17: 32'b11100000000001100110000100000110;
		10'd18: 32'b00010000000100010000001010010001;
		10'd19: 32'b00000000100000010101000010010111;
		10'd20: 32'b00000001000011110000000100010011;
		10'd21: 32'b00000100101000010000000000001101;
		10'd22: 32'b00010100000100010001000100010010;
		10'd23: 32'b01101000000000000000000000111000;
		10'd24: 32'b01000000000010010100000100000010;
		10'd25: 32'b00100000001000010010000100100001;
		10'd26: 32'b00110000001100010010000100010000;
		10'd27: 32'b00000000110100100000000111000111;
		10'd28: 32'b00000011000100100001000100000110;
		10'd29: 32'b00010100000100110001000000100000;
		10'd30: 32'b00010001001000101011000110100110;
		10'd31: 32'b10000000000100001000010000001010;
		10'd32: 32'b10010000110000001001000100010000;
		10'd33: 32'b01000100010000010100001001010000;
		10'd34: 32'b00110000000000011100000100001010;
		10'd35: 32'b00000001000110100000000100010101;
		10'd36: 32'b01000000010100000100001001010010;
		10'd37: 32'b00000000011000000001010001110000;
		10'd38: 32'b00010010000000100001001000000110;
		10'd39: 32'b00100000000010011000010000000010;
		10'd40: 32'b00011000100000010000100100000010;
		10'd41: 32'b00000010000000111110000000001110;
		10'd42: 32'b01000000001100100000000100100110;
		10'd43: 32'b00000000000000010110001100100011;
		10'd44: 32'b00100000000000010010100100010001;
		10'd45: 32'b00010001000100000000001100000010;
		10'd46: 32'b00011000110000010010000001000000;
		10'd47: 32'b11000101000010000100000100100000;
		10'd48: 32'b00000001100100000000000111010000;
		10'd49: 32'b10101000000001001011000000000000;
		10'd50: 32'b01010000000000110000010100000111;
		10'd51: 32'b01000001010100010100000100000101;
		10'd52: 32'b10000100000010101000010100000001;
		10'd53: 32'b00000101000001000000011001010110;
		10'd54: 32'b01010000000101100101000000000110;
		10'd55: 32'b00011000000000010001100100001001;
		10'd56: 32'b00000000100100110000000011010101;
		10'd57: 32'b00100001000001110000000100000001;
		10'd58: 32'b00010001010000010000010001000010;
		10'd59: 32'b10010000000001101001000000000110;
		10'd60: 32'b00100000000001110001000100000110;
		10'd61: 32'b01100000100001000010000010000000;
		10'd62: 32'b01000010010000110100001100010001;
		10'd63: 32'b11110011000110111011110110011001;
		10'd64: 32'b11101111111111101100010101111000;
		10'd65: 32'b11110000110110111011010101111111;
		10'd66: 32'b11111101111001001011000101001101;
		10'd67: 32'b11000011011110110111010101000000;
		10'd68: 32'b01110111111111101100100011010100;
		10'd69: 32'b01010111101010110110100101110000;
		10'd70: 32'b10100111100000111011011101101011;
		10'd71: 32'b10111110011010010101001000011011;
		10'd72: 32'b11010101100110111010110100101011;
		10'd73: 32'b11000101001001110110011101011101;
		10'd74: 32'b11110111000101110011001000001011;
		10'd75: 32'b10000101011000110011011110000010;
		10'd76: 32'b10111100010011011111011110011001;
		10'd77: 32'b10000001010011010001001101011001;
		10'd78: 32'b11110101011101111111001110111111;
		10'd79: 32'b11101010011010111110111101110001;
		10'd80: 32'b01010110000111011110011001101011;
		10'd81: 32'b00001110111010101111110011000110;
		10'd82: 32'b01010001011101000011011000101100;
		10'd83: 32'b11011010111101001101001000110011;
		10'd84: 32'b01100110000010110111110101001001;
		10'd85: 32'b10011010011010100011110011111101;
		10'd86: 32'b11000000001110100011111011100110;
		10'd87: 32'b00101100001011011010101111010101;
		10'd88: 32'b10011101101011111110100111110001;
		10'd89: 32'b01000111010111110011001010100101;
		10'd90: 32'b11111001001111100011001110000111;
		10'd91: 32'b00101101000010010010011001010111;
		10'd92: 32'b01000111111101100000101101101011;
		10'd93: 32'b00110111011111001100111100110011;
		10'd94: 32'b01100010101001000001111101011111;
		10'd95: 32'b01101101010111010010010111001011;
		10'd96: 32'b00011010000101010101000010001001;
		10'd97: 32'b10001111010101011000111010001111;
		10'd98: 32'b10110101101011110101011111000111;
		10'd99: 32'b11000100010010010110110000000101;
		10'd100: 32'b01101110111001010110001000001001;
		10'd101: 32'b11011011010011110000111100001011;
		10'd102: 32'b00111111000001111001000101000001;
		10'd103: 32'b10101111100011100011001010001101;
		10'd104: 32'b11010111110111111110100100111100;
		10'd105: 32'b10011111111101101000011110111010;
		10'd106: 32'b00010011111111100110110010010011;
		10'd107: 32'b00101111110101111000001110111100;
		10'd108: 32'b11111111111101011011111100011100;
		10'd109: 32'b00001011111010101111010101011101;
		10'd110: 32'b01011011111110101100011001101101;
		10'd111: 32'b00111100111011111111011111111010;
		10'd112: 32'b11110101000101100111001101110111;
		10'd113: 32'b00000100010100000111101001110011;
		10'd114: 32'b11110011000111101101111001101111;
		10'd115: 32'b00110110000011111101001011100111;
		10'd116: 32'b11100011111001101110010000111011;
		10'd117: 32'b11011010000111100111001011110111;
		10'd118: 32'b11011001001111101000101011110011;
		10'd119: 32'b00111000010100100011100001010110;
		10'd120: 32'b10010100100010011011010011110010;
		10'd121: 32'b01110110000100100001100000011111;
		10'd122: 32'b10110101010100100001010011111111;
		10'd123: 32'b00111110000000000011101011010010;
		10'd124: 32'b10011100010001011100100100110111;
		10'd125: 32'b10110111011110000100110100010110;
		10'd126: 32'b11111011100100010100110110111111;
		10'd127: 32'b01111011001011001111101110010001;
		10'd128: 32'b11111011111100111110110000100010;
		10'd129: 32'b00100111011111001111001010011101;
		10'd130: 32'b11111111101110101011100111110111;
		10'd131: 32'b01001111001011000100000101111011;
		10'd132: 32'b10011001101101001110110010000010;
		10'd133: 32'b00100100111011000001100011011110;
		10'd134: 32'b11111011111111101111100101111111;
		10'd135: 32'b10111101011100111000100111101000;
		10'd136: 32'b11111101000100111111101000100010;
		10'd137: 32'b11100101110001111010111000001101;
		10'd138: 32'b11111111111111101011100110010101;
		10'd139: 32'b10001111110100101011110001101010;
		10'd140: 32'b00111010101110011000101101111000;
		10'd141: 32'b01111111110001111111111110001101;
		10'd142: 32'b11111111110111100001101110001100;
		10'd143: 32'b00111100011101010100010000110010;
		10'd144: 32'b11100010111011001010100010111111;
		10'd145: 32'b00101100110110101111111001001001;
		10'd146: 32'b11111101111010111100100010101001;
		10'd147: 32'b00100100001011001101111100010011;
		10'd148: 32'b00111000110111011110110011100111;
		10'd149: 32'b10100010010010011111011111010000;
		10'd150: 32'b10111010111010001110100011101011;
		10'd151: 32'b10000101100001010110000110011001;
		10'd152: 32'b11001111111111011110110110001100;
		10'd153: 32'b00111010100011111110010001101010;
		10'd154: 32'b11111001110011011010100110111000;
		10'd155: 32'b10101011111111000110110110011011;
		10'd156: 32'b11111011010100110111000010101000;
		10'd157: 32'b01110001100010001110000011101110;
		10'd158: 32'b11111101111010111100011010011100;
		10'd159: 32'b00110000110101110001100110111001;
		10'd160: 32'b01111110101111100101101001110000;
		10'd161: 32'b11111000100111010001101010011010;
		10'd162: 32'b11110111100101100000011100110100;
		10'd163: 32'b01011111100001101011101101010011;
		10'd164: 32'b11010111111111001000101111101010;
		10'd165: 32'b11101000100100000101111000010101;
		10'd166: 32'b01110001101010000110001111111100;
		10'd167: 32'b10010111110001110011100110011110;
		10'd168: 32'b01100110110011110010110111000111;
		10'd169: 32'b00011100011011100000011010100100;
		10'd170: 32'b10011011100011000010111100010100;
		10'd171: 32'b01001101000001010101111110111111;
		10'd172: 32'b00101100100110001000110110110100;
		10'd173: 32'b00001100011011111001010010001111;
		10'd174: 32'b01010001100111010011111101011100;
		10'd175: 32'b01110101000100010000111101100111;
		10'd176: 32'b11010000000011100011111001111000;
		10'd177: 32'b11010111011111000000111111111111;
		10'd178: 32'b00001110000000000000011111111001;
		10'd179: 32'b11010111000101000000001011011011;
		10'd180: 32'b11000110111001000101111011111010;
		10'd181: 32'b10101110011111000001101110110110;
		10'd182: 32'b10011011101000010011001011111001;
		10'd183: 32'b01110110010000011011000010100110;
		10'd184: 32'b11001110101101110100111011101111;
		10'd185: 32'b11110001101101010000111100111001;
		10'd186: 32'b11110000100001011001110110101110;
		10'd187: 32'b01110010001110011001001011100100;
		10'd188: 32'b00010100111111111111111110110101;
		10'd189: 32'b11110000001110101000011111100110;
		10'd190: 32'b11110111101101100010110110110110;
		10'd191: 32'b01011100010110101001011110011101;
		10'd192: 32'b01001001001100001101010110001101;
		10'd193: 32'b00000111011111010101111001101011;
		10'd194: 32'b11011100000001000011101110100110;
		10'd195: 32'b01000010111100111110111001001111;
		10'd196: 32'b01110100110100000100110000011101;
		10'd197: 32'b10111001011110101011001101110011;
		10'd198: 32'b00111101000011101000000101101100;
		10'd199: 32'b00100010111111010101010101000111;
		10'd200: 32'b00001000011111100101111011000000;
		10'd201: 32'b01110000110001001110110110011101;
		10'd202: 32'b01110101010101000110010001100101;
		10'd203: 32'b01010011110001010101010101010101;
		10'd204: 32'b11101110100110011110000111110001;
		10'd205: 32'b01110011110010010111110100011001;
		10'd206: 32'b01111101101001001110011011100111;
		10'd207: 32'b01111001010010101000010110101000;
		10'd208: 32'b01101111001001011010001011010110;
		10'd209: 32'b01001111000101100001110110101100;
		10'd210: 32'b00010110110110010110110011100000;
		10'd211: 32'b11111010110000111000001111000110;
		10'd212: 32'b01000111101100110011101110111011;
		10'd213: 32'b01001011110100100010100111101001;
		10'd214: 32'b00000001011001100011010001111011;
		10'd215: 32'b10001001111001011110110000111101;
		10'd216: 32'b10100101101001000111000010000110;
		10'd217: 32'b01100111111100101111001110011101;
		10'd218: 32'b00110100001011111010001001010010;
		10'd219: 32'b11010100111111101011011100011101;
		10'd220: 32'b00000101111001010110010111100000;
		10'd221: 32'b01111001011111001111110110111100;
		10'd222: 32'b10000100111101111010010010010110;
		10'd223: 32'b10111011101101111000011100100101;
		10'd224: 32'b10010101010010111101001100111110;
		10'd225: 32'b01111101011111111100100110100010;
		10'd226: 32'b10110001110111101101000110101100;
		10'd227: 32'b10000111100101111111101110000010;
		10'd228: 32'b10011110010010011011100100110110;
		10'd229: 32'b10101011001010010101100110101010;
		10'd230: 32'b11011011111100111101001110110101;
		10'd231: 32'b10100011101110111001110111000110;
		10'd232: 32'b10100101101101000111101100101010;
		10'd233: 32'b11010101111111111111111110111110;
		10'd234: 32'b01100101100011001111000111101111;
		10'd235: 32'b00110101001100100000110010101010;
		10'd236: 32'b11111100101100101001101001101010;
		10'd237: 32'b10101001110100110101111101111100;
		10'd238: 32'b10100000101110000100011111111000;
		10'd239: 32'b10001101111000100111101110111000;
		10'd240: 32'b00001000001000110100111110001011;
		10'd241: 32'b11111101110100000001010111110100;
		10'd242: 32'b10001111101101111010101111000000;
		10'd243: 32'b11001101100010000111101110111011;
		10'd244: 32'b00110010000101111110111111010001;
		10'd245: 32'b11000011101100011111100110101100;
		10'd246: 32'b00111101101000100011110010001010;
		10'd247: 32'b10001011100000110111101010111110;
		10'd248: 32'b11110101101010110000000111101011;
		10'd249: 32'b11110000000011101011011110011101;
		10'd250: 32'b11010011101101111000001011100001;
		10'd251: 32'b10010100010001110001111110001101;
		10'd252: 32'b11111011010101111010000011101011;
		10'd253: 32'b01100101000011010001101111011000;
		10'd254: 32'b01000011111000110001010111111011;
		10'd255: 32'b01000100010111001110010101011010;
		10'd256: 32'b11001101110000001111111111011101;
		10'd257: 32'b11000010010101101110010101010010;
		10'd258: 32'b11001001110000100011010010110011;
		10'd259: 32'b11001011011101011111111111000010;
		10'd260: 32'b11101011100000111111111111011101;
		10'd261: 32'b01010110010101111110110101111110;
		10'd262: 32'b01000101110000100111011111111100;
		10'd263: 32'b00111001101101100001111001101110;
		10'd264: 32'b11111101010101101110110010010011;
		10'd265: 32'b10101010111100100001111100011111;
		10'd266: 32'b01101001011100110110110011011001;
		10'd267: 32'b10111001000101100011111110010110;
		10'd268: 32'b10111101111101110111100010011011;
		10'd269: 32'b10100000010101100111100010110111;
		10'd270: 32'b10111001101101101001110001111111;
		10'd271: 32'b00101111110100110100100101011011;
		10'd272: 32'b01001101111111100110001100101101;
		10'd273: 32'b01100101111011000101010000110010;
		10'd274: 32'b01110111011110101011010111000000;
		10'd275: 32'b01111111110001001101110101111010;
		10'd276: 32'b11111101111010001101100100011000;
		10'd277: 32'b00100011110011101000101011001111;
		10'd278: 32'b01111101111101100111000000000000;
		10'd279: 32'b11011100011110110000111110010010;
		10'd280: 32'b11010101001011011001010111011011;
		10'd281: 32'b10110111101111010100111110110001;
		10'd282: 32'b11100101111100011011111110010000;
		10'd283: 32'b11001101001110110010111011110100;
		10'd284: 32'b11011110101010011000011010010001;
		10'd285: 32'b10011100101011011110100111111000;
		10'd286: 32'b11001111110010011000101010011010;
		10'd287: 32'b01100001011100101110111011111101;
		10'd288: 32'b10111010101100011111011011000101;
		10'd289: 32'b11011101111100001011010110111010;
		10'd290: 32'b11110111111110111010111101001011;
		10'd291: 32'b11111111110100111010100111110000;
		10'd292: 32'b10110101111100111011011010000011;
		10'd293: 32'b11111110110101111011110111000111;
		10'd294: 32'b11110101011110110010001111111101;
		10'd295: 32'b00111110011011001011110111101011;
		10'd296: 32'b11110110011110101111011110111110;
		10'd297: 32'b01011010110001101000011101010011;
		10'd298: 32'b11000011000011001001011010110100;
		10'd299: 32'b00010010100011000100110110001110;
		10'd300: 32'b11011010101011110010000000101000;
		10'd301: 32'b10000101111011111111100100000010;
		10'd302: 32'b11001111110011100101110111110011;
		10'd303: 32'b10101100111011110110111000110010;
		10'd304: 32'b10010101000010111001001111100111;
		10'd305: 32'b00111011111101111111101110010101;
		10'd306: 32'b00101101010000110110001001001111;
		10'd307: 32'b01101100110011100110111100010110;
		10'd308: 32'b10101101111001101000111100000100;
		10'd309: 32'b01010101011111111110101000001000;
		10'd310: 32'b01101100111001110011101000111111;
		10'd311: 32'b01100011011001011111010110110000;
		10'd312: 32'b01000001001000110111110010101111;
		10'd313: 32'b11001101101101110001110011011110;
		10'd314: 32'b10011000010000101011100010001010;
		10'd315: 32'b11110110010001011101110110000110;
		10'd316: 32'b01110000111101011001010010001011;
		10'd317: 32'b11100011111101111011000111000010;
		10'd318: 32'b11111010011010011000010011011010;
		10'd319: 32'b10010111111000110101010111011001;
		10'd320: 32'b11001011101001111111011100001000;
		10'd321: 32'b10011111111010111111001100111111;
		10'd322: 32'b00011111111110111101011100100001;
		10'd323: 32'b11110110111001010011100010000011;
		10'd324: 32'b00011111001100111111111101110100;
		10'd325: 32'b11001100111110110101000101111111;
		10'd326: 32'b11010111111110111111010010101001;
		10'd327: 32'b10101111111010111001111010110111;
		10'd328: 32'b11100101011011111010011101001111;
		10'd329: 32'b10101111001110100010000011111110;
		10'd330: 32'b00101001110010011100011111111101;
		10'd331: 32'b10100011101000011001111011011101;
		10'd332: 32'b11100100111111111010111101100011;
		10'd333: 32'b00111011101111000111010111001111;
		10'd334: 32'b11110101011101011001010111011001;
		10'd335: 32'b10111011010101011001111001011001;
		10'd336: 32'b10100100010001000000101101111100;
		10'd337: 32'b10011111011000000110110000001011;
		10'd338: 32'b11001100111000000000010110111111;
		10'd339: 32'b11110011010110010101111001001011;
		10'd340: 32'b10001001111110000111111101011011;
		10'd341: 32'b10111010110011000011011101101111;
		10'd342: 32'b11001111101000010010110100101011;
		10'd343: 32'b11011111110110001110101111101111;
		10'd344: 32'b10111011010101110101000010111100;
		10'd345: 32'b10001011110111110110111010100111;
		10'd346: 32'b10100001011000010100110111100111;
		10'd347: 32'b11001101110011111100111100011001;
		10'd348: 32'b10100000111111011100010110110100;
		10'd349: 32'b11100111110110110110010100001111;
		10'd350: 32'b10001001011010000100011000000101;
		10'd351: 32'b11101101001111001010101010101101;
		10'd352: 32'b00101111101101110111000011110011;
		10'd353: 32'b11011001111010010010111110101001;
		10'd354: 32'b11110010110000010010111011101100;
		10'd355: 32'b00101110111011010010101100101011;
		10'd356: 32'b00111011101001010000011011001001;
		10'd357: 32'b00101010010110110001001110101011;
		10'd358: 32'b10000110100001111010111000111101;
		10'd359: 32'b11101001000010101011011110101100;
		10'd360: 32'b11100010000111101110011010110000;
		10'd361: 32'b01001110000110011000010110011100;
		10'd362: 32'b01111111100001001111011000111101;
		10'd363: 32'b11011001001100001010011110111101;
		10'd364: 32'b11000111000110101001011100101010;
		10'd365: 32'b11001101111000111110000010101110;
		10'd366: 32'b11000111100111001110011001100100;
		10'd367: 32'b10101001111011101110001111111001;
		10'd368: 32'b01011110111100111101011011000100;
		10'd369: 32'b01111111101011010111001100001000;
		10'd370: 32'b10001011100101001001011111101111;
		10'd371: 32'b10100001101010111010101110101101;
		10'd372: 32'b11101110111101100001000101100101;
		10'd373: 32'b11111001010101000111110010100001;
		10'd374: 32'b11000111011000000001101111111111;
		10'd375: 32'b11001001100000110111011011111111;
		10'd376: 32'b00111101101100100101011011011111;
		10'd377: 32'b01011101101110100011100111111111;
		10'd378: 32'b00111001100011011011111011111111;
		10'd379: 32'b01011000111010000101000011111111;
		10'd380: 32'b01111001101010100101110101011011;
		10'd381: 32'b00111101101101110010010011010111;
		10'd382: 32'b00111101101101010011011011111110;
		10'd383: 32'b10011111010011100001010100110000;
		10'd384: 32'b11011111010111011111001001011110;
		10'd385: 32'b10101111010110101011110111111000;
		10'd386: 32'b11010110001010110111101100001010;
		10'd387: 32'b10011101011000001011111111110011;
		10'd388: 32'b10011111011100101001110101010001;
		10'd389: 32'b10100101100010011010010110111010;
		10'd390: 32'b11110011011010010101110000010111;
		10'd391: 32'b01101100010100001111110011011101;
		10'd392: 32'b01111111101110110110011110001011;
		10'd393: 32'b01100011110100001110010101111110;
		10'd394: 32'b11111001111100000101101111011010;
		10'd395: 32'b01111011100011101000111010011100;
		10'd396: 32'b10111100110111110101011111011110;
		10'd397: 32'b11101110111100101111011110011010;
		10'd398: 32'b00100011111111101100011010011010;
		10'd399: 32'b01010111111001110001010000110111;
		10'd400: 32'b10100100010000001111111110110110;
		10'd401: 32'b11010011010001100000110000111001;
		10'd402: 32'b01110110111100001000100111111101;
		10'd403: 32'b11000111000000100100011001111101;
		10'd404: 32'b10010110111000110111010011110111;
		10'd405: 32'b11110111011110110010111001111110;
		10'd406: 32'b11010111111010101110011101111111;
		10'd407: 32'b10011000100110110011111111110101;
		10'd408: 32'b00110110101111111111011111100101;
		10'd409: 32'b00111110101111111101110111000110;
		10'd410: 32'b01111011111100111001111010010010;
		10'd411: 32'b01111100100100101100111101010101;
		10'd412: 32'b10111110111110101011110111001101;
		10'd413: 32'b00011111010111111001000111100101;
		10'd414: 32'b10010100111100111001111111000101;
		10'd415: 32'b00111110011100001111111101001010;
		10'd416: 32'b10101010001111100001011011111001;
		10'd417: 32'b10111011011100100010011011000101;
		10'd418: 32'b11101101111111100111111111011101;
		10'd419: 32'b11101010101001010111111101010100;
		10'd420: 32'b01110000101111100101010011110111;
		10'd421: 32'b10111011101101100010011101000010;
		10'd422: 32'b10111100111011100101110001011111;
		10'd423: 32'b10111011111000101110000011010100;
		10'd424: 32'b10111011100001110010010100010110;
		10'd425: 32'b11111000010010011000100110110110;
		10'd426: 32'b01101101101011010011111110011010;
		10'd427: 32'b10011001101111110000010011000001;
		10'd428: 32'b10111001101011110000100100111000;
		10'd429: 32'b10111001101100011000010110000110;
		10'd430: 32'b11000101101111111001111100011111;
		10'd431: 32'b11110111001100110111001100101001;
		10'd432: 32'b10100111110000000111011011000110;
		10'd433: 32'b00100101101101000110010111010010;
		10'd434: 32'b11101111011100010100111110101101;
		10'd435: 32'b11110000100101000110001100000100;
		10'd436: 32'b00110010111001111111111110000011;
		10'd437: 32'b01110001010100001111101010101001;
		10'd438: 32'b11001010110000100111111001111000;
		10'd439: 32'b11010111111111011100110010001010;
		10'd440: 32'b10011001001111100011011001011111;
		10'd441: 32'b01001101001111101001101001110110;
		10'd442: 32'b10011101010110100011011100110110;
		10'd443: 32'b11011110001110111000110110110010;
		10'd444: 32'b10010100000110101101011000010111;
		10'd445: 32'b00011101111110111001100010100010;
		10'd446: 32'b11011100100110010011011111100110;
		10'd447: 32'b10001000111110011001101010100111;
		10'd448: 32'b10011111101010011111101111011111;
		10'd449: 32'b01111111101000010111111110001101;
		10'd450: 32'b00110010100110111110111010011011;
		10'd451: 32'b10111001110011111111111111110001;
		10'd452: 32'b10111011111100100111011111111111;
		10'd453: 32'b00010010011100010111101010000111;
		10'd454: 32'b11110001111010011111111000001010;
		10'd455: 32'b00001111101000001110100101110111;
		10'd456: 32'b00001010011100000111100100011001;
		10'd457: 32'b01000111111101101101100110111011;
		10'd458: 32'b11001010110110101100100110111000;
		10'd459: 32'b00101111101000011011101110110100;
		10'd460: 32'b10111010011111111000101100111001;
		10'd461: 32'b11101010001001000011110101110111;
		10'd462: 32'b00011011000000001011100000010000;
		10'd463: 32'b11100001000011000110011100001010;
		10'd464: 32'b00110100011110001100100001000000;
		10'd465: 32'b00110000101010001000100010111001;
		10'd466: 32'b10110011111011101110110011011011;
		10'd467: 32'b00100100110010101011011001111111;
		10'd468: 32'b10000111110010001110110000001010;
		10'd469: 32'b00100100111110000100111000001010;
		10'd470: 32'b11110101011011010000100111101011;
		10'd471: 32'b00111110000001100110111100110000;
		10'd472: 32'b01111101101110100110110000110001;
		10'd473: 32'b01100011010010000010100010111001;
		10'd474: 32'b00011001100101000110111010100111;
		10'd475: 32'b01010011001100111110101000100100;
		10'd476: 32'b01001110010001110111011001111101;
		10'd477: 32'b01111001010001101010111011110000;
		10'd478: 32'b00101011010001000110111000111101;
		10'd479: 32'b10111010000010001110011010000000;
		10'd480: 32'b01110010011101001011100101110001;
		10'd481: 32'b11101110001001001110111111000110;
		10'd482: 32'b01100100010100111110001011000011;
		10'd483: 32'b01111010011011010110111010111101;
		10'd484: 32'b10100000111111001101101001110110;
		10'd485: 32'b11111000100001101100101011011010;
		10'd486: 32'b00100110011101001010110100001101;
		10'd487: 32'b10111101001110011000111000101101;
		10'd488: 32'b00100110111010001000011101101110;
		10'd489: 32'b11110001011011111010101000001111;
		10'd490: 32'b00010000111011111001110001100011;
		10'd491: 32'b10101101111000111000011101101111;
		10'd492: 32'b10101110111001101000101000110110;
		10'd493: 32'b00100010111111001000101100111101;
		10'd494: 32'b10101100111000011001110010000011;
		10'd495: 32'b00010101101111010010011101111001;
		10'd496: 32'b11110010011100100101001000101110;
		10'd497: 32'b00110111001010110000011100011100;
		10'd498: 32'b01111010111110101101001000111101;
		10'd499: 32'b00010101011011010111101110011001;
		10'd500: 32'b10110110001001001111000001111100;
		10'd501: 32'b01100110110010111000010010001000;
		10'd502: 32'b10111111001110100110101010111100;
		10'd503: 32'b01001111100101111000111010111111;
		10'd504: 32'b01011111101011111010011111111111;
		10'd505: 32'b11000011101001111101110000010011;
		10'd506: 32'b10100011011111111101000110101011;
		10'd507: 32'b11001110000000110100110001010011;
		10'd508: 32'b00111100110110100000111100100001;
		10'd509: 32'b11100010010100011011110000010001;
		10'd510: 32'b10111110001101110110000100101101;
		10'd511: 32'b01101101011101100010011101111011;
		10'd512: 32'b01000101001000110000111011110010;
		10'd513: 32'b01111011110101010010111110101111;
		10'd514: 32'b11010111101101111101101110111010;
		10'd515: 32'b11101101001001010011110110101110;
		10'd516: 32'b01011001101101110010100110110111;
		10'd517: 32'b01101001100100010100111111010010;
		10'd518: 32'b11110111011101110011111010110011;
		10'd519: 32'b11111101101011001010100101011111;
		10'd520: 32'b10111001100111010001111100101100;
		10'd521: 32'b10101100001011100000011011111001;
		10'd522: 32'b11111101101111101100111110111111;
		10'd523: 32'b00011110111010011110101101100101;
		10'd524: 32'b01011110010111000011110010011110;
		10'd525: 32'b01011001101001111110111100111011;
		10'd526: 32'b11110101101111001100100101100101;
		10'd527: 32'b00110011000011000101010000010110;
		10'd528: 32'b11110011011000101001100111111010;
		10'd529: 32'b11110001000001110111101001011110;
		10'd530: 32'b10100011001101000001100100000010;
		10'd531: 32'b11100011100010011001001101110010;
		10'd532: 32'b01111101011001100101101111010010;
		10'd533: 32'b01111101001101110011010011111111;
		10'd534: 32'b11101001001111111001100111010110;
		10'd535: 32'b11101101110000101111111000111110;
		10'd536: 32'b01110101011101001111100010011110;
		10'd537: 32'b10111110111111101011100100100000;
		10'd538: 32'b00100110101011011010110010110101;
		10'd539: 32'b11101001100111001011111110100111;
		10'd540: 32'b10111110011001000110101011110100;
		10'd541: 32'b10110110011001101110111010010001;
		10'd542: 32'b10011000011110001111111011101111;
		10'd543: 32'b01110000111010011100001101000110;
		10'd544: 32'b00001011110101010110101111111101;
		10'd545: 32'b11110011110100011010010011110111;
		10'd546: 32'b00100111110101000001101001110100;
		10'd547: 32'b00111000111011000000100010000000;
		10'd548: 32'b00011110110101001010100001000100;
		10'd549: 32'b00010101101101000011111110010011;
		10'd550: 32'b00100011110001111101101001001101;
		10'd551: 32'b01101011011111010100111000111000;
		10'd552: 32'b10101011111100111111011110000111;
		10'd553: 32'b00101001111110111010110100111100;
		10'd554: 32'b11100000010110001010110110100011;
		10'd555: 32'b11011001001100110101110001111101;
		10'd556: 32'b00101111101111111110101111001101;
		10'd557: 32'b01100011110111001110111001111101;
		10'd558: 32'b11011011001100110100110111001110;
		10'd559: 32'b11111000110110010111100011011100;
		10'd560: 32'b11101010011101100100001011010010;
		10'd561: 32'b01011011111100111000000111101011;
		10'd562: 32'b00101000101101111101101011101101;
		10'd563: 32'b01111001111111111011100111001101;
		10'd564: 32'b01101000101100100110001011100100;
		10'd565: 32'b00001111011000010001000001001111;
		10'd566: 32'b00101100101011111000100011110110;
		10'd567: 32'b00100111011011000000010000110100;
		10'd568: 32'b01111011100011110001111111101001;
		10'd569: 32'b10111111110010111101110110010100;
		10'd570: 32'b01101001011000010001111111010110;
		10'd571: 32'b10110111111111100100000010100100;
		10'd572: 32'b00111011010010001001010111110111;
		10'd573: 32'b00111101110011111111011111001100;
		10'd574: 32'b01111010110000010101111011010100;
	endcase;
	return out;
endfunction
function Bit#(32) get_output_page5(UInt#(10) counter);
	Bit#(32) out = case(counter)
		10'd0: 32'b01000100100011010100010110001000;
		10'd1: 32'b01110000000101000001010000110100;
		10'd2: 32'b00001100011001000000100001100110;
		10'd3: 32'b00010011000000110000001101110010;
		10'd4: 32'b00000101001001000100000101100100;
		10'd5: 32'b10000000010100010000000000010100;
		10'd6: 32'b01010001000010100101000101011011;
		10'd7: 32'b01000010010000110001001101000110;
		10'd8: 32'b10000101110000000010000101000010;
		10'd9: 32'b01000101011001110100010001010101;
		10'd10: 32'b00010001100001110000000110000110;
		10'd11: 32'b00010001000100010001000000011011;
		10'd12: 32'b00000000010110000100010101100100;
		10'd13: 32'b00000000101000100000000000110101;
		10'd14: 32'b00000100001101110000010000100100;
		10'd15: 32'b01000000010000000111000111000000;
		10'd16: 32'b00011010010001110001110000000111;
		10'd17: 32'b11100000000001100110000100100110;
		10'd18: 32'b00010000000100110000001010010001;
		10'd19: 32'b10000000100000010101000010010111;
		10'd20: 32'b00010001000011110000000100011011;
		10'd21: 32'b00000110101000010000000000001101;
		10'd22: 32'b00010101000100110001000100010010;
		10'd23: 32'b01101100000000000000000000111010;
		10'd24: 32'b01000001001010010100000100100011;
		10'd25: 32'b00110000001100010010000100100001;
		10'd26: 32'b00110000001100010010000100010100;
		10'd27: 32'b00000010110101100000000111000111;
		10'd28: 32'b00000011010100100001000100000110;
		10'd29: 32'b00011100000100110001000000100000;
		10'd30: 32'b10110001101000101011000110110110;
		10'd31: 32'b10000000000101001000010000001010;
		10'd32: 32'b10010000110000001001000111010000;
		10'd33: 32'b01000101010000010100011001010000;
		10'd34: 32'b00110000000000111100010100001010;
		10'd35: 32'b00000001000110100010000100010101;
		10'd36: 32'b01000000110100000100001001010010;
		10'd37: 32'b00000100011000010001010001110000;
		10'd38: 32'b01010010000000100001001000000110;
		10'd39: 32'b00100000100010111000010010000011;
		10'd40: 32'b00111000100000010000100110000010;
		10'd41: 32'b00000010000000111111001000001110;
		10'd42: 32'b01001000001100100010000100101110;
		10'd43: 32'b00100000000000010110001100100011;
		10'd44: 32'b00101001000010010010100100010001;
		10'd45: 32'b00010011000100000100001100000010;
		10'd46: 32'b00011000110000110011000001000000;
		10'd47: 32'b11100101001010000100000100100001;
		10'd48: 32'b00010001110100000100000111010000;
		10'd49: 32'b10101000000001001011100100000000;
		10'd50: 32'b01010001000100110001010100000111;
		10'd51: 32'b01000001010100010100001101000101;
		10'd52: 32'b11000100000010101000010100001001;
		10'd53: 32'b00100101010001000000011001010110;
		10'd54: 32'b01010010000101100101000000010110;
		10'd55: 32'b00011000000010010001100100001101;
		10'd56: 32'b00000000100100111000000011010101;
		10'd57: 32'b00100001000001110000001100010001;
		10'd58: 32'b00010101010000110000010001000010;
		10'd59: 32'b10010000000001101011001000100110;
		10'd60: 32'b00100001000001110001000100000110;
		10'd61: 32'b01100000100101000110000010000000;
		10'd62: 32'b01010010010100110100001101010011;
		10'd63: 32'b11110011110110111011110110011001;
		10'd64: 32'b11101111111111101100010101111100;
		10'd65: 32'b11110001110111111011110101111111;
		10'd66: 32'b11111101111101111111001101001101;
		10'd67: 32'b11010111011110110111010111001000;
		10'd68: 32'b11110111111111111111110111110101;
		10'd69: 32'b01010111101110110110110101110010;
		10'd70: 32'b11100111101010111011011111101111;
		10'd71: 32'b10111110111010010101011001011011;
		10'd72: 32'b11010101101111111110110100111011;
		10'd73: 32'b11000101011001111110011101011101;
		10'd74: 32'b11110111000101110011001000011011;
		10'd75: 32'b10000111011000110111011110000011;
		10'd76: 32'b10111100110011011111011111011011;
		10'd77: 32'b10000101011011010001001101011001;
		10'd78: 32'b11110111011101111111001110111111;
		10'd79: 32'b11101110011010111110111101110001;
		10'd80: 32'b01110110000111011110011001101011;
		10'd81: 32'b00001110111011101111110011000110;
		10'd82: 32'b11010011011101100011011000101100;
		10'd83: 32'b11011010111101011101001000110011;
		10'd84: 32'b01100110000110110111110111001001;
		10'd85: 32'b10111010011010100011110011111101;
		10'd86: 32'b11000001001110100011111011100110;
		10'd87: 32'b00101100011011011010101111010101;
		10'd88: 32'b10011101101011111110101111111001;
		10'd89: 32'b11000111011111110011001010100101;
		10'd90: 32'b11111001001111101011001110000111;
		10'd91: 32'b10101101001011110010011001010111;
		10'd92: 32'b01000111111111100001101101101011;
		10'd93: 32'b00110111011111001100111100111011;
		10'd94: 32'b01100011101101010001111101011111;
		10'd95: 32'b01101101010111010010110111001011;
		10'd96: 32'b00111010000101010101000011001001;
		10'd97: 32'b10011111010111011000111011001111;
		10'd98: 32'b10111101111011110101011111001111;
		10'd99: 32'b11000100010011010110111000001101;
		10'd100: 32'b01111110111001010110011011001001;
		10'd101: 32'b11011011010011110000111110011111;
		10'd102: 32'b00111111100001111101000101000001;
		10'd103: 32'b10111111110111100011001010111101;
		10'd104: 32'b11010111110111111111110100111100;
		10'd105: 32'b10011111111111101000011111111010;
		10'd106: 32'b00010011111111100110110110010111;
		10'd107: 32'b10101111110101111000011110111100;
		10'd108: 32'b11111111111101111111111100011110;
		10'd109: 32'b10011011111010101111110101011101;
		10'd110: 32'b01011011111110101100011001101111;
		10'd111: 32'b00111100111011111111011111111010;
		10'd112: 32'b11110101001101100111111101110111;
		10'd113: 32'b00000100010100001111101001110011;
		10'd114: 32'b11110011000111101101111011101111;
		10'd115: 32'b00110110000011111111001011101111;
		10'd116: 32'b11100011111001111110010000111011;
		10'd117: 32'b11011010001111100111001011110111;
		10'd118: 32'b11111011001111101100101111110111;
		10'd119: 32'b00111010010100100011100001010110;
		10'd120: 32'b10010100100010011111110011110011;
		10'd121: 32'b01110110000100110001101000011111;
		10'd122: 32'b10110101110100100011010011111111;
		10'd123: 32'b01111110000100000011101011010010;
		10'd124: 32'b10011100010011011100100110110111;
		10'd125: 32'b11110111011111100100110100010111;
		10'd126: 32'b11111111100100010100110110111111;
		10'd127: 32'b01111011001111101111101111010001;
		10'd128: 32'b11111011111101111110110000100010;
		10'd129: 32'b00100111011111001111101010011101;
		10'd130: 32'b11111111101110101111110111110111;
		10'd131: 32'b01001111111011000101000101111011;
		10'd132: 32'b11111001101101001110110010000010;
		10'd133: 32'b10110100111011000011100011011110;
		10'd134: 32'b11111011111111101111100111111111;
		10'd135: 32'b10111111111100111101100111101000;
		10'd136: 32'b11111111000100111111101100100010;
		10'd137: 32'b11100101110011111011111000001101;
		10'd138: 32'b11111111111111101011101110010101;
		10'd139: 32'b10011111110100111011111001101010;
		10'd140: 32'b01111010101110011000101101111000;
		10'd141: 32'b11111111110001111111111110001101;
		10'd142: 32'b11111111110111101001101110001100;
		10'd143: 32'b01111100011101010100010000110010;
		10'd144: 32'b11100110111011001110101010111111;
		10'd145: 32'b00101110110110101111111001001001;
		10'd146: 32'b11111101111010111100100110101001;
		10'd147: 32'b00100100001011001101111101010011;
		10'd148: 32'b00111000110111011110110011100111;
		10'd149: 32'b10100010010011011111011111010000;
		10'd150: 32'b10111010111011001110110011101011;
		10'd151: 32'b10001111100011010110000110011001;
		10'd152: 32'b11001111111111011110110110101101;
		10'd153: 32'b00111011101011111110010011101010;
		10'd154: 32'b11111001110011011110100110111000;
		10'd155: 32'b10101011111111000110110110011011;
		10'd156: 32'b11111011110110110111000110101100;
		10'd157: 32'b01111001100011001110010111111110;
		10'd158: 32'b11111101111111111100011010011100;
		10'd159: 32'b01110000110111110001100111111001;
		10'd160: 32'b01111110101111110101101001110000;
		10'd161: 32'b11111000100111010001101110011010;
		10'd162: 32'b11110111100101100011011110110100;
		10'd163: 32'b01011111100001101011101101011011;
		10'd164: 32'b11011111111111001000111111101010;
		10'd165: 32'b11111010100100100111111010010101;
		10'd166: 32'b01111011101011000110011111111100;
		10'd167: 32'b10010111110001110011101110011110;
		10'd168: 32'b01100110110011110110111111110111;
		10'd169: 32'b00111100111011101000011010111100;
		10'd170: 32'b10011011100011101010111100010100;
		10'd171: 32'b01001111010001110101111110111111;
		10'd172: 32'b00101100110110001000111110110100;
		10'd173: 32'b00001101011111111001110010101111;
		10'd174: 32'b11010011100111010011111101011100;
		10'd175: 32'b11110101001100010000111111110111;
		10'd176: 32'b11010100010111100011111011111000;
		10'd177: 32'b11010111011111000010111111111111;
		10'd178: 32'b00011111001100000000111111111011;
		10'd179: 32'b11110111000101000000011011011011;
		10'd180: 32'b11000110111001001101111011111010;
		10'd181: 32'b11111110111111000101111110110110;
		10'd182: 32'b10011111101000010011101011111001;
		10'd183: 32'b01110110011100011011001010100110;
		10'd184: 32'b11011110101111110100111011101111;
		10'd185: 32'b11110001101101110000111110111001;
		10'd186: 32'b11110010101001011001110110101111;
		10'd187: 32'b01110010001110011001001011101101;
		10'd188: 32'b00010110111111111111111110110101;
		10'd189: 32'b11110110001110101001111111100111;
		10'd190: 32'b11110111101101100010110111110110;
		10'd191: 32'b01011101010110101011011110011101;
		10'd192: 32'b11011001011110001111010110001101;
		10'd193: 32'b00000111011111111111111001101011;
		10'd194: 32'b11011100010001000011111110100110;
		10'd195: 32'b01000010111100111110111001001111;
		10'd196: 32'b01110100111100000100110100011101;
		10'd197: 32'b10111001011110101011001101110011;
		10'd198: 32'b00111101000011101010001101101100;
		10'd199: 32'b00110010111111010101010101010111;
		10'd200: 32'b01101100011111111101111111100100;
		10'd201: 32'b01110000110001011110111110011101;
		10'd202: 32'b01111101010111010111010001100101;
		10'd203: 32'b01010011110001010101110101011101;
		10'd204: 32'b11101110110110111110000111110001;
		10'd205: 32'b01110011110011010111110100011001;
		10'd206: 32'b01111101101101001110011011101111;
		10'd207: 32'b11111001010010111000010110101000;
		10'd208: 32'b01111111001001111011001111111110;
		10'd209: 32'b01001111000101110101110110101100;
		10'd210: 32'b00010110111110010110111111100001;
		10'd211: 32'b11111011110010111000101111100110;
		10'd212: 32'b01000111101100111111101110111011;
		10'd213: 32'b01001011110101100010100111111001;
		10'd214: 32'b00010011011101110011010001111111;
		10'd215: 32'b11011001111001011111110011111101;
		10'd216: 32'b10100111101001001111001010101110;
		10'd217: 32'b01100111111100101111001110011101;
		10'd218: 32'b10110100011111111110001101010110;
		10'd219: 32'b11111100111111101111111100011101;
		10'd220: 32'b10000101111001010111010111110100;
		10'd221: 32'b11111001011111101111110110111100;
		10'd222: 32'b11000100111101111010010011010110;
		10'd223: 32'b10111011111101111000111100100101;
		10'd224: 32'b10010111010010111101101100111110;
		10'd225: 32'b01111101011111111100101110100010;
		10'd226: 32'b11110001111111111101001111101100;
		10'd227: 32'b10110111101101111111111110010010;
		10'd228: 32'b10011110010110011011100100111110;
		10'd229: 32'b10101011001011011101100110101010;
		10'd230: 32'b11111111111100111101001110110101;
		10'd231: 32'b10100011101110111001110111010110;
		10'd232: 32'b10100101111101100111101100111010;
		10'd233: 32'b11010111111111111111111110111110;
		10'd234: 32'b01100101110011001111110111101111;
		10'd235: 32'b00110101101100100010110010101010;
		10'd236: 32'b11111110101100101001101101111110;
		10'd237: 32'b10111001111100110111111101111110;
		10'd238: 32'b10100000101110100100011111111010;
		10'd239: 32'b10001101111000100111101110111000;
		10'd240: 32'b00101000001000110100111110001011;
		10'd241: 32'b11111101110100000001010111110100;
		10'd242: 32'b10111111101101111010111111000100;
		10'd243: 32'b11001111100010000111101110111011;
		10'd244: 32'b00110010100101111110111111010001;
		10'd245: 32'b11000011101100011111100110101100;
		10'd246: 32'b10111101111000100011110010001110;
		10'd247: 32'b11011011100100110111101010111110;
		10'd248: 32'b11110101101110110000000111101011;
		10'd249: 32'b11110100000111101011011110011101;
		10'd250: 32'b11010011101101111000001111100011;
		10'd251: 32'b10010101010001110001111111011101;
		10'd252: 32'b11111011010101111011000011101011;
		10'd253: 32'b01100101000011011001111111011000;
		10'd254: 32'b11100011111000110001010111111011;
		10'd255: 32'b01000110010111011111010101011110;
		10'd256: 32'b11001101110000101111111111011101;
		10'd257: 32'b11000010010101101110111101010010;
		10'd258: 32'b11001101110010110011010010110111;
		10'd259: 32'b11001011111101111111111111010110;
		10'd260: 32'b11101011101000111111111111011101;
		10'd261: 32'b01010110010111111110111101111111;
		10'd262: 32'b01000111110000100111011111111101;
		10'd263: 32'b00111001111111101111111101101111;
		10'd264: 32'b11111101010101101110110110011011;
		10'd265: 32'b10101111111100110001111100011111;
		10'd266: 32'b01111011011100111111110011011001;
		10'd267: 32'b11111101000101100011111110110110;
		10'd268: 32'b10111101111111110111110010011011;
		10'd269: 32'b10101000010101100111100010111111;
		10'd270: 32'b10111001101101101011110001111111;
		10'd271: 32'b00101111110101110110100101011011;
		10'd272: 32'b01001101111111101111001110101101;
		10'd273: 32'b01100101111011001101010000110010;
		10'd274: 32'b01111111111110101011010111000000;
		10'd275: 32'b01111111111001001101110101111011;
		10'd276: 32'b11111101111010001111110100011100;
		10'd277: 32'b00101111111111101010101011001111;
		10'd278: 32'b01111101111111110111000111000000;
		10'd279: 32'b11011100111110110000111110010010;
		10'd280: 32'b11010101001011011001011111111111;
		10'd281: 32'b10110111101111011100111110110101;
		10'd282: 32'b11100101111100011011111110010010;
		10'd283: 32'b11001101001110111010111011110100;
		10'd284: 32'b11011110101010011000011010010001;
		10'd285: 32'b11011100101011011110110111111000;
		10'd286: 32'b11101111111011111011111010011011;
		10'd287: 32'b11110001111100101110111111111101;
		10'd288: 32'b11111111101100111111011011000101;
		10'd289: 32'b11011101111100011011110111111111;
		10'd290: 32'b11110111111110111010111101101011;
		10'd291: 32'b11111111111100111010101111110100;
		10'd292: 32'b10110101111101111011011011000011;
		10'd293: 32'b11111110110101111011110111010111;
		10'd294: 32'b11110101111111111011001111111101;
		10'd295: 32'b00111111011011001011110111101111;
		10'd296: 32'b11110110011110101111011110111110;
		10'd297: 32'b01011110110011101000011111010011;
		10'd298: 32'b11010011000111101011011110110100;
		10'd299: 32'b00010010100011000100110110011110;
		10'd300: 32'b11011010111111110010000000101000;
		10'd301: 32'b10110101111011111111100101011010;
		10'd302: 32'b11001111110011100101110111111011;
		10'd303: 32'b10101101111011110110111000110011;
		10'd304: 32'b10010101000010111001001111100111;
		10'd305: 32'b00111011111101111111101110011101;
		10'd306: 32'b00111101010000110111001001001111;
		10'd307: 32'b01101100110011100111111100010111;
		10'd308: 32'b10101101111001101000111100001100;
		10'd309: 32'b01011101011111111111101100001100;
		10'd310: 32'b01101100111001111011111000111111;
		10'd311: 32'b01100111011001011111010110110010;
		10'd312: 32'b01000011001000111111110010101111;
		10'd313: 32'b11001111101101110001111011111110;
		10'd314: 32'b11011000110000111011110010001011;
		10'd315: 32'b11110110010011011101110110000110;
		10'd316: 32'b01110000111111011011110010001011;
		10'd317: 32'b11100011111101111011000111100010;
		10'd318: 32'b11111010011010111000010011011010;
		10'd319: 32'b10010111111000110101010111011001;
		10'd320: 32'b11011011101001111111111100101000;
		10'd321: 32'b10011111111010111111001101111111;
		10'd322: 32'b11111111111110111101111100100001;
		10'd323: 32'b11110110111001110011100111101011;
		10'd324: 32'b00011111011100111111111101110100;
		10'd325: 32'b11001100111111110101000101111111;
		10'd326: 32'b11010111111110111111010110101001;
		10'd327: 32'b10101111111010111001111110110111;
		10'd328: 32'b11100101111011111010011101101111;
		10'd329: 32'b10101111011110101011010111111110;
		10'd330: 32'b01101101111010011100011111111101;
		10'd331: 32'b10100011111000011001111111011101;
		10'd332: 32'b11100100111111111111111101100011;
		10'd333: 32'b00111111101111100111111111001111;
		10'd334: 32'b11110111111101011001010111011111;
		10'd335: 32'b10111111010101111101111001011001;
		10'd336: 32'b10100101010011010000101111111100;
		10'd337: 32'b10011111011010010110110000001011;
		10'd338: 32'b11001100111000000000010110111111;
		10'd339: 32'b11110011010110011101111011001011;
		10'd340: 32'b11011101111110010111111101011011;
		10'd341: 32'b10111010110011000011011101101111;
		10'd342: 32'b11001111111000010010110100101011;
		10'd343: 32'b11011111110110011110101111101111;
		10'd344: 32'b10111011010111111101000110111101;
		10'd345: 32'b10001011110111110110111010101111;
		10'd346: 32'b10100001011010010100111111100111;
		10'd347: 32'b11001111110111111100111100111111;
		10'd348: 32'b10100010111111111100010110111100;
		10'd349: 32'b11100111110110110110111100001111;
		10'd350: 32'b10001001011010000100011000100101;
		10'd351: 32'b11101101101111001010101010101111;
		10'd352: 32'b00101111101101111111001011111011;
		10'd353: 32'b11011111111110010010111110101001;
		10'd354: 32'b11110010110000010010111011101100;
		10'd355: 32'b00101111111011010010101100101011;
		10'd356: 32'b00111011101011010000011011101001;
		10'd357: 32'b00101011110110110001001110101011;
		10'd358: 32'b10000110101011111010111010111101;
		10'd359: 32'b11101011011110101011011110111101;
		10'd360: 32'b11100110000111101110011110110000;
		10'd361: 32'b01001111000110111010010110111100;
		10'd362: 32'b01111111101001011111111010111101;
		10'd363: 32'b11011001001100001010011110111101;
		10'd364: 32'b11000111000111101001011100101010;
		10'd365: 32'b11001101111000111110001010101110;
		10'd366: 32'b11001111100111001111011001110110;
		10'd367: 32'b10111011111011101110001111111011;
		10'd368: 32'b01011111111100111101011011000100;
		10'd369: 32'b01111111101111010111001100101010;
		10'd370: 32'b10001011100101001001011111101111;
		10'd371: 32'b10100001101010111011101110101101;
		10'd372: 32'b11101111111101101001000101101101;
		10'd373: 32'b11111001010101000111110010100001;
		10'd374: 32'b11001111011000000101101111111111;
		10'd375: 32'b11001101100000110111011111111111;
		10'd376: 32'b00111101101100110101011011011111;
		10'd377: 32'b01011101101111110111110111111111;
		10'd378: 32'b00111101101011011011111011111111;
		10'd379: 32'b01011000111010010101010011111111;
		10'd380: 32'b01111101101110100101110111011011;
		10'd381: 32'b00111101101111110011011011110111;
		10'd382: 32'b01111101101101011011011011111110;
		10'd383: 32'b10111111010011100001010100110000;
		10'd384: 32'b11011111010111111111011001011110;
		10'd385: 32'b10101111010110101011110111111010;
		10'd386: 32'b11010110101010110111101110001010;
		10'd387: 32'b10011111011000011011111111110011;
		10'd388: 32'b10011111011110111001110101010001;
		10'd389: 32'b10110101110110011010011110111010;
		10'd390: 32'b11110111011110010101110000011111;
		10'd391: 32'b01101100110100001111110011011101;
		10'd392: 32'b01111111111110110111011111011011;
		10'd393: 32'b01100011111100001111010101111110;
		10'd394: 32'b11111101111110000101101111011011;
		10'd395: 32'b01111011110011101110111010011100;
		10'd396: 32'b11111100110111110101011111011110;
		10'd397: 32'b11101110111100101111011110011010;
		10'd398: 32'b00100011111111101100011010111010;
		10'd399: 32'b01010111111001111001010000110111;
		10'd400: 32'b10100110010100001111111110110110;
		10'd401: 32'b11010011010001100001110000111001;
		10'd402: 32'b01110111111100101000100111111111;
		10'd403: 32'b11000111000001100100011101111101;
		10'd404: 32'b10010110111000110111010011110111;
		10'd405: 32'b11110111011110110011111001111110;
		10'd406: 32'b11010111111110101110011101111111;
		10'd407: 32'b10011000100110110011111111110101;
		10'd408: 32'b00110110101111111111011111100101;
		10'd409: 32'b00111110101111111101110111110110;
		10'd410: 32'b01111111111101111101111111011010;
		10'd411: 32'b01111100100110101101111101110101;
		10'd412: 32'b10111110111110101111110111011101;
		10'd413: 32'b00011111110111111001011111100101;
		10'd414: 32'b10011100111100111001111111000101;
		10'd415: 32'b01111110011100011111111101001011;
		10'd416: 32'b10101010001111101101011011111001;
		10'd417: 32'b11111011111100100011011011000101;
		10'd418: 32'b11101101111111100111111111011111;
		10'd419: 32'b11101010101001110111111101010110;
		10'd420: 32'b01110100101111101101010011110111;
		10'd421: 32'b10111011111101110010011101100010;
		10'd422: 32'b10111100111011100111110101011111;
		10'd423: 32'b10111011111000101110000011010100;
		10'd424: 32'b10111011100001110011010100010110;
		10'd425: 32'b11111000010010011000100110110110;
		10'd426: 32'b01101101101011010011111110011010;
		10'd427: 32'b10011001101111110000010111000001;
		10'd428: 32'b10111011101011110000100100111010;
		10'd429: 32'b10111001101100111001010110100110;
		10'd430: 32'b11001111101111111001111100011111;
		10'd431: 32'b11110111101100110111111100101001;
		10'd432: 32'b10100111110000000111011011001110;
		10'd433: 32'b01100101111101010110011111010010;
		10'd434: 32'b11101111111100010100111110101111;
		10'd435: 32'b11110000100101100110001100100100;
		10'd436: 32'b11110010111001111111111110000011;
		10'd437: 32'b01110011010100001111101010101001;
		10'd438: 32'b11111010110000100111111011111000;
		10'd439: 32'b11010111111111111100110010111010;
		10'd440: 32'b10111001001111100011011101011111;
		10'd441: 32'b11001101001111101001101001110110;
		10'd442: 32'b10011111011110100011011101110110;
		10'd443: 32'b11011110001110111000110110110010;
		10'd444: 32'b10010101000110101101111000110111;
		10'd445: 32'b00011101111110111001100010111010;
		10'd446: 32'b11011100100110010011011111100110;
		10'd447: 32'b10111010111110111101111010101111;
		10'd448: 32'b10011111101010011111101111011111;
		10'd449: 32'b01111111111000010111111110001111;
		10'd450: 32'b00111010101110111110111010011011;
		10'd451: 32'b11111001111011111111111111110001;
		10'd452: 32'b10111011111100100111011111111111;
		10'd453: 32'b00010010011110010111111010001111;
		10'd454: 32'b11110001111010011111111110001010;
		10'd455: 32'b00001111101000001110100101111111;
		10'd456: 32'b00001010011100110111100100011001;
		10'd457: 32'b01101111111101101101100110111111;
		10'd458: 32'b11001011110110111100100110111011;
		10'd459: 32'b00101111101000011011101110110100;
		10'd460: 32'b10111011011111111000101101111011;
		10'd461: 32'b11111010011001100011110101110111;
		10'd462: 32'b10111011110000001011100000010001;
		10'd463: 32'b11100001000011000110011100001010;
		10'd464: 32'b00110100011110011100100001011001;
		10'd465: 32'b00110000101110001000100010111011;
		10'd466: 32'b10110011111011101110110011011011;
		10'd467: 32'b00100100110010101011111001111111;
		10'd468: 32'b10000111110010101110111000001010;
		10'd469: 32'b00100110111110000110111001001010;
		10'd470: 32'b11110111011011010100100111101011;
		10'd471: 32'b00111111001001100110111100110000;
		10'd472: 32'b01111101101111100110110001110001;
		10'd473: 32'b01100011011010000010100111111001;
		10'd474: 32'b01111101100101000111111010100111;
		10'd475: 32'b01010011011100111110101000100100;
		10'd476: 32'b01101110010001110111111001111101;
		10'd477: 32'b01111001010001101010111011110001;
		10'd478: 32'b00111011010001010110111000111101;
		10'd479: 32'b11111010100111001110011010100100;
		10'd480: 32'b01110010111101001011101101110001;
		10'd481: 32'b11111110001001001110111111000111;
		10'd482: 32'b01111100010100111110101111010011;
		10'd483: 32'b11111010011011110110111010111101;
		10'd484: 32'b10100000111111001101101001110110;
		10'd485: 32'b11111000111011101100101011011010;
		10'd486: 32'b00101110011101011110110110001101;
		10'd487: 32'b11111101011110011000111000101101;
		10'd488: 32'b00100110111011011000111101111110;
		10'd489: 32'b11110001011011111010111000001111;
		10'd490: 32'b01010100111011111001111001100111;
		10'd491: 32'b10101101111000111000111101101111;
		10'd492: 32'b10111110111001101000111001110110;
		10'd493: 32'b10101011111111001000101100111101;
		10'd494: 32'b10101100111001011001110010010011;
		10'd495: 32'b00010101101111010011111101111001;
		10'd496: 32'b11111010011100100101001000101110;
		10'd497: 32'b00110111011011110000011100011100;
		10'd498: 32'b01111110111110101101101000111101;
		10'd499: 32'b00010101011011110111101110011001;
		10'd500: 32'b10110110001011001111000001111100;
		10'd501: 32'b01110110111010111000010010001000;
		10'd502: 32'b10111111001110100110101010111100;
		10'd503: 32'b01101111100101111001111010111111;
		10'd504: 32'b01011111101011111011011111111111;
		10'd505: 32'b11010011101001111101110000010011;
		10'd506: 32'b10100011111111111101000110101011;
		10'd507: 32'b11001110000000110100110001010011;
		10'd508: 32'b00111100111111111101111100110001;
		10'd509: 32'b11100110010100011011110000110011;
		10'd510: 32'b11111110001111111110110100101111;
		10'd511: 32'b11101101011101100010011111111111;
		10'd512: 32'b01010101101100110000111011110010;
		10'd513: 32'b01111111110101010010111110101111;
		10'd514: 32'b11011111101111111101101110111110;
		10'd515: 32'b11101111001101011011110111111110;
		10'd516: 32'b01011001101111110010111110110111;
		10'd517: 32'b01111001110100010100111111011111;
		10'd518: 32'b11110111111101110111111010110111;
		10'd519: 32'b11111101101011011010111101011111;
		10'd520: 32'b10111001100111110001111100101100;
		10'd521: 32'b10101100101011100001111011111001;
		10'd522: 32'b11111101101111101101111110111111;
		10'd523: 32'b00011110111010011110101101100101;
		10'd524: 32'b11011110010111000011110111011110;
		10'd525: 32'b01011001101001111110111101111011;
		10'd526: 32'b11111101101111001100101101110101;
		10'd527: 32'b01110011100011000111010000010110;
		10'd528: 32'b11111011011000101001100111111010;
		10'd529: 32'b11110001000001110111111101111110;
		10'd530: 32'b10110011101101010001100110000010;
		10'd531: 32'b11110011100010011001011101110010;
		10'd532: 32'b01111101011001100101101111111010;
		10'd533: 32'b11111101001111110011010011111111;
		10'd534: 32'b11101001001111111001100111010110;
		10'd535: 32'b11101101111011101111111000111110;
		10'd536: 32'b01110101111101101111110010111110;
		10'd537: 32'b10111110111111101011100100100000;
		10'd538: 32'b01100110101011011010110011110111;
		10'd539: 32'b11101001100111001111111110100111;
		10'd540: 32'b10111110011001011110101011111100;
		10'd541: 32'b11111110011001101110111110010011;
		10'd542: 32'b10111010111110001111111111111111;
		10'd543: 32'b01110000111010011100001111010110;
		10'd544: 32'b00011011110101111110101111111101;
		10'd545: 32'b11111011110100011010010011111111;
		10'd546: 32'b00100111110101100001101001110100;
		10'd547: 32'b00111000111011000100110010000110;
		10'd548: 32'b00011111110101001010100101000101;
		10'd549: 32'b00010101111101000111111110011011;
		10'd550: 32'b00110011110001111101111001001101;
		10'd551: 32'b01101011011111110100111101111000;
		10'd552: 32'b10101011111100111111111110100111;
		10'd553: 32'b00101001111110111010110100111100;
		10'd554: 32'b11100011110110001010110111100011;
		10'd555: 32'b11011001101100110101111001111101;
		10'd556: 32'b11101111111111111110101111001101;
		10'd557: 32'b01101011110111101110111001111101;
		10'd558: 32'b11011011011101111110110111101110;
		10'd559: 32'b11111000110111010111100011011100;
		10'd560: 32'b11101010111101100111001011010110;
		10'd561: 32'b01111011111100111001000111101111;
		10'd562: 32'b00101010101111111101101011101101;
		10'd563: 32'b11111001111111111011100111001101;
		10'd564: 32'b01111010101100101110001011111100;
		10'd565: 32'b00001111111000111011000011101111;
		10'd566: 32'b00101100101111111001100011110110;
		10'd567: 32'b00100111111111000010010000110100;
		10'd568: 32'b01111111100011110001111111101101;
		10'd569: 32'b10111111110011111101110111110100;
		10'd570: 32'b01101101011000010001111111010110;
		10'd571: 32'b10110111111111100100000010100100;
		10'd572: 32'b00111011010010001001110111110111;
		10'd573: 32'b00111101110011111111011111001101;
		10'd574: 32'b01111010110111011101111011010101;
	endcase;
	return out;
endfunction
function Bit#(32) get_output_page6(UInt#(10) counter);
	Bit#(32) out = case(counter)
		10'd0: 32'b01000100100011110100010110001000;
		10'd1: 32'b01110000000111000001010000110100;
		10'd2: 32'b00001110011001000000100001100110;
		10'd3: 32'b00010111000100110001011101110011;
		10'd4: 32'b00000101001101010100000101100100;
		10'd5: 32'b10000000110101011000000010010100;
		10'd6: 32'b01110001001010110101001101011011;
		10'd7: 32'b01000010010000111001001101000110;
		10'd8: 32'b10000101110000000010000101000010;
		10'd9: 32'b01010101011001110100010011010101;
		10'd10: 32'b00010001100001110000000110010111;
		10'd11: 32'b00010001000100011001000100011011;
		10'd12: 32'b00000000010110000100010101110100;
		10'd13: 32'b00100000101000100000000010110101;
		10'd14: 32'b00000100001101110000010100100101;
		10'd15: 32'b01000000110000000111000111000000;
		10'd16: 32'b00011110010001110001110001000111;
		10'd17: 32'b11100000100001100110000110100110;
		10'd18: 32'b11010000000100110000001010010001;
		10'd19: 32'b10010000100000010101000010010111;
		10'd20: 32'b00010001010011110000001100011011;
		10'd21: 32'b00001110101010010000000000001101;
		10'd22: 32'b00011101000100110001000100010010;
		10'd23: 32'b01101100000000000000010000111010;
		10'd24: 32'b01000001001010010100000100101011;
		10'd25: 32'b00110000001100010010000100100001;
		10'd26: 32'b00110100001101010010010100010101;
		10'd27: 32'b00100010110101100000000111000111;
		10'd28: 32'b00000111010100100001010101000110;
		10'd29: 32'b00011100001110110001000000100000;
		10'd30: 32'b10110011101100101011000110110111;
		10'd31: 32'b10100000000101001000010000001010;
		10'd32: 32'b11010001110100001101000111010000;
		10'd33: 32'b01000101010000010100111001010000;
		10'd34: 32'b00110100000000111100010100001110;
		10'd35: 32'b00000001001110100010000100011101;
		10'd36: 32'b01000000110100000100001001010110;
		10'd37: 32'b00000100011000010001010001110011;
		10'd38: 32'b01010011000000100101001000000110;
		10'd39: 32'b00100001100010111100010010000011;
		10'd40: 32'b00111001100000010000100110000110;
		10'd41: 32'b00000010000000111111001100011110;
		10'd42: 32'b01101000001100110110000100101111;
		10'd43: 32'b10100000000000010110001100101011;
		10'd44: 32'b00101001010010010010100100010101;
		10'd45: 32'b01010011000100000100001100000011;
		10'd46: 32'b00011000110001110011010001010000;
		10'd47: 32'b11100101001010000100000101100001;
		10'd48: 32'b01010001110101000100000111010000;
		10'd49: 32'b10101000000001001011100110000000;
		10'd50: 32'b01010101001100110101010100100111;
		10'd51: 32'b01000001010100010110001101010101;
		10'd52: 32'b11000101000010101100010100001001;
		10'd53: 32'b00100101010101000000011001010110;
		10'd54: 32'b01010011000101100101000001010110;
		10'd55: 32'b00011000000011010001100100011101;
		10'd56: 32'b00001000100100111000001011010101;
		10'd57: 32'b00100001000001110001001100110011;
		10'd58: 32'b00010101010000110000010001000110;
		10'd59: 32'b11010010000001101011001000100110;
		10'd60: 32'b00100001000101110001000100000110;
		10'd61: 32'b01100000100101001110100010001000;
		10'd62: 32'b01010110010100110101001101010111;
		10'd63: 32'b11110011110110111111110111011001;
		10'd64: 32'b11101111111111101101010101111100;
		10'd65: 32'b11110001110111111111110101111111;
		10'd66: 32'b11111101111101111111001101001101;
		10'd67: 32'b11010111011110110111010111101010;
		10'd68: 32'b11110111111111111111110111111101;
		10'd69: 32'b01010111111111110110110101110010;
		10'd70: 32'b11100111101011111011011111101111;
		10'd71: 32'b10111110111011010101011001011011;
		10'd72: 32'b11110101111111111111111100111011;
		10'd73: 32'b11000101011001111111011101011101;
		10'd74: 32'b11110111000111110011001000011011;
		10'd75: 32'b10000111011000110111011110000011;
		10'd76: 32'b10111110110111011111011111011011;
		10'd77: 32'b10000101011011010001011111011101;
		10'd78: 32'b11110111011101111111001110111111;
		10'd79: 32'b11101110011010111111111101110001;
		10'd80: 32'b01110110000111011110011001101011;
		10'd81: 32'b00001110111011101111110011000110;
		10'd82: 32'b11011011011101100011011000101100;
		10'd83: 32'b11011010111101011101001000110011;
		10'd84: 32'b01100110000110110111110111101001;
		10'd85: 32'b10111010011010100011110011111101;
		10'd86: 32'b11000001001110110011111011100110;
		10'd87: 32'b00111100011011011010101111010101;
		10'd88: 32'b10011101101011111110101111111001;
		10'd89: 32'b11000111011111110011001010100101;
		10'd90: 32'b11111001001111101011001110000111;
		10'd91: 32'b10101101001011111010011001010111;
		10'd92: 32'b01000111111111100001101111101011;
		10'd93: 32'b00110111011111001100111100111011;
		10'd94: 32'b01100011101101010001111111011111;
		10'd95: 32'b01101101010111010010110111001011;
		10'd96: 32'b01111010000101010101000011001001;
		10'd97: 32'b10011111010111011000111011011111;
		10'd98: 32'b10111101111011110101011111001111;
		10'd99: 32'b11000100010011110110111010001101;
		10'd100: 32'b01111111111001010110011011001001;
		10'd101: 32'b11011011010011110000111110011111;
		10'd102: 32'b00111111100001111101010101000111;
		10'd103: 32'b10111111110111100011001010111101;
		10'd104: 32'b11010111110111111111110100111100;
		10'd105: 32'b10011111111111101000011111111010;
		10'd106: 32'b00010011111111100110110110010111;
		10'd107: 32'b10101111110101111000011110111100;
		10'd108: 32'b11111111111101111111111100011110;
		10'd109: 32'b10011011111111101111111101011101;
		10'd110: 32'b01011011111111101100011001101111;
		10'd111: 32'b00111100111011111111011111111010;
		10'd112: 32'b11110101101101100111111101110111;
		10'd113: 32'b00100100010100101111101001111011;
		10'd114: 32'b11110011000111101101111011101111;
		10'd115: 32'b00111110001011111111001011101111;
		10'd116: 32'b11100011111001111110011000111011;
		10'd117: 32'b11011010011111100111001011110111;
		10'd118: 32'b11111111001111101100101111110111;
		10'd119: 32'b00111110110100100011100001010110;
		10'd120: 32'b10110100100010011111110011110111;
		10'd121: 32'b01110110001100110001101000011111;
		10'd122: 32'b10110101110100100011010011111111;
		10'd123: 32'b01111110000100000011101011010010;
		10'd124: 32'b10011100010011011100100110111111;
		10'd125: 32'b11110111011111100100110110010111;
		10'd126: 32'b11111111100101010100110110111111;
		10'd127: 32'b01111011001111101111101111010001;
		10'd128: 32'b11111011111111111110110000100010;
		10'd129: 32'b00100111111111001111101010011111;
		10'd130: 32'b11111111101110101111110111110111;
		10'd131: 32'b11001111111011001101000111111011;
		10'd132: 32'b11111001101101001110111010000010;
		10'd133: 32'b10110100111011010011100011011110;
		10'd134: 32'b11111011111111101111100111111111;
		10'd135: 32'b10111111111100111101101111101000;
		10'd136: 32'b11111111100110111111101100101010;
		10'd137: 32'b11101111110011111011111000001101;
		10'd138: 32'b11111111111111101011101110010101;
		10'd139: 32'b10011111110100111011111001101010;
		10'd140: 32'b11111010101110011000101101111000;
		10'd141: 32'b11111111110001111111111110001101;
		10'd142: 32'b11111111110111101001101110001100;
		10'd143: 32'b01111100011101010100010000110010;
		10'd144: 32'b11100110111011001110101010111111;
		10'd145: 32'b00101110110110101111111001001001;
		10'd146: 32'b11111101111010111100100110101001;
		10'd147: 32'b00100100001011001101111101010011;
		10'd148: 32'b00111000111111011110110011100111;
		10'd149: 32'b10100110010011011111011111010000;
		10'd150: 32'b10111010111011001110110011101011;
		10'd151: 32'b10001111100011010110010110011001;
		10'd152: 32'b11001111111111011111110110101101;
		10'd153: 32'b00111011101011111110010011101010;
		10'd154: 32'b11111001110011011110100110111000;
		10'd155: 32'b10101011111111000110111110011011;
		10'd156: 32'b11111011110110110111100110101100;
		10'd157: 32'b11111001100011001110010111111110;
		10'd158: 32'b11111101111111111100011010011100;
		10'd159: 32'b01110000110111110001100111111001;
		10'd160: 32'b01111110101111110111111001110000;
		10'd161: 32'b11111000100111010001101111011010;
		10'd162: 32'b11110111100101100011011111110100;
		10'd163: 32'b01011111100111101011101101111011;
		10'd164: 32'b11011111111111001000111111101110;
		10'd165: 32'b11111010100101100111111010010101;
		10'd166: 32'b01111011101111000111111111111100;
		10'd167: 32'b10010111110011110011101110011110;
		10'd168: 32'b01100110110011110110111111110111;
		10'd169: 32'b00111100111011111001111010111100;
		10'd170: 32'b10011011100011101011111100010100;
		10'd171: 32'b01001111011001110111111110111111;
		10'd172: 32'b00101100110110001000111110110100;
		10'd173: 32'b00001101011111111001110010111111;
		10'd174: 32'b11010011100111010011111101011100;
		10'd175: 32'b11110101001110010000111111110111;
		10'd176: 32'b11010100010111100011111011111000;
		10'd177: 32'b11010111011111000010111111111111;
		10'd178: 32'b00011111001100000000111111111011;
		10'd179: 32'b11110111000101000000011011011011;
		10'd180: 32'b11010110111001001101111011111010;
		10'd181: 32'b11111111111111100101111110111110;
		10'd182: 32'b10011111101000010011111011111011;
		10'd183: 32'b01110111011100011011001010110110;
		10'd184: 32'b11011110101111110100111111111111;
		10'd185: 32'b11110001101101110000111110111001;
		10'd186: 32'b11110010101101011001110110101111;
		10'd187: 32'b01110010001110011001001011111101;
		10'd188: 32'b00010110111111111111111110110101;
		10'd189: 32'b11110110001111101001111111100111;
		10'd190: 32'b11110111101101100010110111110110;
		10'd191: 32'b01011101010110101011011110111101;
		10'd192: 32'b11011001011110001111010110001111;
		10'd193: 32'b00010111011111111111111101101011;
		10'd194: 32'b11111100010101100011111110100110;
		10'd195: 32'b01010010111100111110111001001111;
		10'd196: 32'b01110100111101001101110100011101;
		10'd197: 32'b10111011011110101011001101110011;
		10'd198: 32'b00111101011011111010001101101100;
		10'd199: 32'b01110010111111010101010101010111;
		10'd200: 32'b01101100011111111101111111100111;
		10'd201: 32'b01110000110011011110111110011101;
		10'd202: 32'b01111101010111010111010101100101;
		10'd203: 32'b01011011110001010101110101011101;
		10'd204: 32'b11101110110110111111000111110001;
		10'd205: 32'b01111011110011010111110100011001;
		10'd206: 32'b01111101101101001110011011101111;
		10'd207: 32'b11111001010010111000010110101000;
		10'd208: 32'b01111111001001111011001111111110;
		10'd209: 32'b11011111001101110101110111101100;
		10'd210: 32'b00010110111110111110111111100001;
		10'd211: 32'b11111011110010111000101111100110;
		10'd212: 32'b01000111101100111111101110111011;
		10'd213: 32'b01001011110101110010100111111001;
		10'd214: 32'b00010011011101110011010111111111;
		10'd215: 32'b11111101111001011111110011111101;
		10'd216: 32'b10100111111001001111011010111110;
		10'd217: 32'b01100111111100101111001110011101;
		10'd218: 32'b10110100111111111110001101010110;
		10'd219: 32'b11111100111111101111111100011101;
		10'd220: 32'b10000101111001011111010111111101;
		10'd221: 32'b11111011011111101111110110111100;
		10'd222: 32'b11100100111101111010010011110111;
		10'd223: 32'b10111011111101111001111100100101;
		10'd224: 32'b10010111010010111101101101111110;
		10'd225: 32'b01111101011111111100101111100010;
		10'd226: 32'b11110001111111111101001111101100;
		10'd227: 32'b11110111101101111111111110010010;
		10'd228: 32'b10011110010110011011101100111110;
		10'd229: 32'b10111011001011111101110110101010;
		10'd230: 32'b11111111111100111101001110110101;
		10'd231: 32'b10100011101110111001110111011110;
		10'd232: 32'b10100101111101100111101110111010;
		10'd233: 32'b11010111111111111111111110111110;
		10'd234: 32'b01100101110011001111110111101111;
		10'd235: 32'b00110101101100100010110010101010;
		10'd236: 32'b11111111101100101001101101111110;
		10'd237: 32'b10111001111100110111111101111110;
		10'd238: 32'b11100000101110100100011111111011;
		10'd239: 32'b10001101111000110111101110111001;
		10'd240: 32'b10111000001000110100111110001011;
		10'd241: 32'b11111101110100000101010111111100;
		10'd242: 32'b10111111101101111010111111001100;
		10'd243: 32'b11001111100010000111101110111011;
		10'd244: 32'b00110010100101111110111111110001;
		10'd245: 32'b11101011101100011111100111101100;
		10'd246: 32'b10111101111000100011111011001110;
		10'd247: 32'b11011011100100110111101010111110;
		10'd248: 32'b11110101101110110001000111101011;
		10'd249: 32'b11110100000111101011011110011101;
		10'd250: 32'b11010011101101111000001111100011;
		10'd251: 32'b11010111110001110011111111011101;
		10'd252: 32'b11111011010101111111000011101011;
		10'd253: 32'b01100101000011111001111111011000;
		10'd254: 32'b11100011111001110001010111111011;
		10'd255: 32'b01101110011111011111011101011111;
		10'd256: 32'b11001101110000101111111111011101;
		10'd257: 32'b11000010010111111111111101010110;
		10'd258: 32'b11111111110010110011110010110111;
		10'd259: 32'b11001011111101111111111111010110;
		10'd260: 32'b11101011101000111111111111111101;
		10'd261: 32'b11010110010111111110111101111111;
		10'd262: 32'b01000111110001110111011111111101;
		10'd263: 32'b00111001111111101111111111101111;
		10'd264: 32'b11111101010101101110110110011011;
		10'd265: 32'b10101111111100110001111100011111;
		10'd266: 32'b11111011011100111111110011011001;
		10'd267: 32'b11111101000101100011111110110110;
		10'd268: 32'b11111101111111110111110010011011;
		10'd269: 32'b10101000010101100111100010111111;
		10'd270: 32'b10111001101101101011110001111111;
		10'd271: 32'b00101111110101110110100101011011;
		10'd272: 32'b01001101111111101111001110101101;
		10'd273: 32'b01100111111011001101111000110010;
		10'd274: 32'b01111111111110101011010111000000;
		10'd275: 32'b01111111111001001101110101111011;
		10'd276: 32'b11111101111010001111111100011100;
		10'd277: 32'b00101111111111101110101011001111;
		10'd278: 32'b01111101111111110111000111000000;
		10'd279: 32'b11011100111111110000111110010010;
		10'd280: 32'b11010101001011011001011111111111;
		10'd281: 32'b11110111101111011100111110110101;
		10'd282: 32'b11100101111110011011111110110011;
		10'd283: 32'b11001101101110111010111011111100;
		10'd284: 32'b11011110101010011000011110010011;
		10'd285: 32'b11011101101011011110110111111000;
		10'd286: 32'b11101111111011111011111010011011;
		10'd287: 32'b11110001111100101110111111111101;
		10'd288: 32'b11111111111100111111011011000101;
		10'd289: 32'b11011111111100111011110111111111;
		10'd290: 32'b11110111111111111010111111101011;
		10'd291: 32'b11111111111100111010101111110100;
		10'd292: 32'b11110101111111111011011011000011;
		10'd293: 32'b11111110111101111011110111010111;
		10'd294: 32'b11110101111111111011011111111101;
		10'd295: 32'b00111111111011001011110111101111;
		10'd296: 32'b11110110011110101111011110111110;
		10'd297: 32'b01011110110011101100111111010011;
		10'd298: 32'b11010111000111101011011110110100;
		10'd299: 32'b00010010100011000100110111011110;
		10'd300: 32'b11011010111111110010100000101000;
		10'd301: 32'b10110101111011111111100101011010;
		10'd302: 32'b11001111110011100101110111111011;
		10'd303: 32'b10101101111011110110111000110111;
		10'd304: 32'b10010101000110111001001111100111;
		10'd305: 32'b00111011111101111111101110011101;
		10'd306: 32'b00111101010000110111101001001111;
		10'd307: 32'b01101100110011100111111100010111;
		10'd308: 32'b10101101111001101000111100001101;
		10'd309: 32'b01011101011111111111101100001101;
		10'd310: 32'b01101100111001111011111000111111;
		10'd311: 32'b01100111011001011111010110110010;
		10'd312: 32'b01000011011000111111110010101111;
		10'd313: 32'b11001111101101110001111011111110;
		10'd314: 32'b11011000110000111011110110001011;
		10'd315: 32'b11110110010011011111110110000110;
		10'd316: 32'b01110000111111011011110010001011;
		10'd317: 32'b11100011111101111011010111100010;
		10'd318: 32'b11111010011010111000110011011011;
		10'd319: 32'b10010111111000111101010111011001;
		10'd320: 32'b11011011101001111111111100101000;
		10'd321: 32'b10011111111010111111001101111111;
		10'd322: 32'b11111111111110111101111100100001;
		10'd323: 32'b11110110111001110011100111101011;
		10'd324: 32'b00011111111100111111111101110100;
		10'd325: 32'b11001100111111110101000101111111;
		10'd326: 32'b11010111111110111111010110101001;
		10'd327: 32'b10101111111010111001111110110111;
		10'd328: 32'b11100101111011111010011101101111;
		10'd329: 32'b10101111011110101011011111111110;
		10'd330: 32'b01101101111010011100011111111101;
		10'd331: 32'b10100011111010111001111111011101;
		10'd332: 32'b11100100111111111111111101100111;
		10'd333: 32'b00111111111111100111111111001111;
		10'd334: 32'b11110111111101011001011111011111;
		10'd335: 32'b10111111010101111101111001011001;
		10'd336: 32'b10100111010011010000101111111100;
		10'd337: 32'b10011111011010011110111100001011;
		10'd338: 32'b11001100111000000000110110111111;
		10'd339: 32'b11111011010110011101111011001011;
		10'd340: 32'b11011101111111010111111101011011;
		10'd341: 32'b10111010110011000011011101111111;
		10'd342: 32'b11011111111000010010110100111011;
		10'd343: 32'b11011111110110011110101111101111;
		10'd344: 32'b10111011010111111111000110111101;
		10'd345: 32'b10001011111111111110111010101111;
		10'd346: 32'b10100011011011011100111111100111;
		10'd347: 32'b11001111110111111100111100111111;
		10'd348: 32'b10100010111111111100010111111100;
		10'd349: 32'b11100111110110110110111100001111;
		10'd350: 32'b10001001011010000100011000100101;
		10'd351: 32'b11101101101111011010101010101111;
		10'd352: 32'b00101111101101111111101011111011;
		10'd353: 32'b11111111111110010010111110101001;
		10'd354: 32'b11110010110000010010111011101101;
		10'd355: 32'b00101111111011010010101100101011;
		10'd356: 32'b00111011101011010000011011101001;
		10'd357: 32'b00101011110110110001001110101011;
		10'd358: 32'b10000110101011111010111010111101;
		10'd359: 32'b11101011111110101011011110111101;
		10'd360: 32'b11100111000111111111011110110000;
		10'd361: 32'b01001111100110111010011110111101;
		10'd362: 32'b01111111101101011111111010111101;
		10'd363: 32'b11011001001100001010011110111101;
		10'd364: 32'b11000111000111101001111100111010;
		10'd365: 32'b11001101111000111110001110101110;
		10'd366: 32'b11001111100111001111011001110110;
		10'd367: 32'b10111011111011101111001111111011;
		10'd368: 32'b01011111111100111101011011000100;
		10'd369: 32'b01111111101111010111101100101011;
		10'd370: 32'b10001011100101011001011111101111;
		10'd371: 32'b10100101101010111011101111101101;
		10'd372: 32'b11101111111101101001000101101101;
		10'd373: 32'b11111001010101000111111010100001;
		10'd374: 32'b11001111011000000101101111111111;
		10'd375: 32'b11011101100000110111011111111111;
		10'd376: 32'b00111101111100110101011011011111;
		10'd377: 32'b01011101101111110111110111111111;
		10'd378: 32'b00111101111011011011111011111111;
		10'd379: 32'b01011101111011010101010011111111;
		10'd380: 32'b01111101101110100101110111011111;
		10'd381: 32'b00111101101111110011011111110111;
		10'd382: 32'b01111101101101011111011011111110;
		10'd383: 32'b10111111011011100011010101110000;
		10'd384: 32'b11011111010111111111011001011110;
		10'd385: 32'b10101111110110101011111111111010;
		10'd386: 32'b11010110101010110111101110001010;
		10'd387: 32'b10011111011000011011111111110011;
		10'd388: 32'b10011111011111111001110101010111;
		10'd389: 32'b10110101110110011010011110111010;
		10'd390: 32'b11110111011110011101111000011111;
		10'd391: 32'b01101100110110001111110011011101;
		10'd392: 32'b01111111111110110111011111011011;
		10'd393: 32'b01100011111100001111010101111110;
		10'd394: 32'b11111101111110000101111111011011;
		10'd395: 32'b01111011111111101110111010011100;
		10'd396: 32'b11111100110111110111011111011111;
		10'd397: 32'b11101110111100101111011110011011;
		10'd398: 32'b00100011111111101100011110111010;
		10'd399: 32'b11011111111001111001010000111111;
		10'd400: 32'b10100110010100001111111110110110;
		10'd401: 32'b11010011011101100001110000111001;
		10'd402: 32'b01110111111100101000100111111111;
		10'd403: 32'b11010111000101100100011101111101;
		10'd404: 32'b10010110111000110111110011110111;
		10'd405: 32'b11110111011110110011111001111110;
		10'd406: 32'b11010111111110111110011111111111;
		10'd407: 32'b10111000100110110011111111110101;
		10'd408: 32'b00110110101111111111011111100101;
		10'd409: 32'b00111110101111111101110111110110;
		10'd410: 32'b01111111111101111101111111011110;
		10'd411: 32'b01111101100110111101111101110101;
		10'd412: 32'b10111110111110111111110111011101;
		10'd413: 32'b00111111110111111001011111100101;
		10'd414: 32'b10011100111101111001111111000101;
		10'd415: 32'b01111110011100011111111101001011;
		10'd416: 32'b10101010001111101101011011111001;
		10'd417: 32'b11111011111101100011011011001111;
		10'd418: 32'b11101101111111100111111111011111;
		10'd419: 32'b11101010101101110111111101010110;
		10'd420: 32'b01111100101111101101010011110111;
		10'd421: 32'b11111111111101110011011101100010;
		10'd422: 32'b10111100111111100111111101011111;
		10'd423: 32'b10111011111000101110000011010100;
		10'd424: 32'b10111011100001110011010100011110;
		10'd425: 32'b11111001110010011000100110110110;
		10'd426: 32'b01101101101011010011111110011010;
		10'd427: 32'b10011001101111110000010111001001;
		10'd428: 32'b10111011111011110000100100111010;
		10'd429: 32'b10111001101100111001010110110110;
		10'd430: 32'b11101111101111111001111110011111;
		10'd431: 32'b11110111101100110111111100101101;
		10'd432: 32'b11100111110000010111011011001110;
		10'd433: 32'b01100101111101010110011111010110;
		10'd434: 32'b11101111111100010100111110111111;
		10'd435: 32'b11110100100101100110001100111100;
		10'd436: 32'b11110011111001111111111111001011;
		10'd437: 32'b01110011010100001111101110101101;
		10'd438: 32'b11111010110000100111111011111000;
		10'd439: 32'b11010111111111111100110010111010;
		10'd440: 32'b10111001001111100011011101011111;
		10'd441: 32'b11001101001111101001101001110110;
		10'd442: 32'b10011111011110100011011101110110;
		10'd443: 32'b11011110001110111000110110110010;
		10'd444: 32'b10011101000110101101111010110111;
		10'd445: 32'b00011101111110111001100010111010;
		10'd446: 32'b11011100100110010011011111100110;
		10'd447: 32'b10111010111110111101111011101111;
		10'd448: 32'b10011111111010011111101111011111;
		10'd449: 32'b01111111111000010111111110001111;
		10'd450: 32'b10111010101110111110111011011011;
		10'd451: 32'b11111001111011111111111111110001;
		10'd452: 32'b10111111111100100111011111111111;
		10'd453: 32'b00010110011110010111111010001111;
		10'd454: 32'b11110001111010011111111110001010;
		10'd455: 32'b00001111101000001110100101111111;
		10'd456: 32'b00001010011101111111101100011001;
		10'd457: 32'b01101111111101101111100110111111;
		10'd458: 32'b11001011110110111101100110111011;
		10'd459: 32'b00101111111000011011101111111100;
		10'd460: 32'b10111011011111111001101101111011;
		10'd461: 32'b11111010011001100011110101110111;
		10'd462: 32'b10111011110100001011100000011001;
		10'd463: 32'b11100001000111000110011100001010;
		10'd464: 32'b00111100111110011100100001011001;
		10'd465: 32'b00110000101110001010100010111011;
		10'd466: 32'b10110111111011101110110011011011;
		10'd467: 32'b10100100110010101011111001111111;
		10'd468: 32'b10001111110010101110111000011010;
		10'd469: 32'b00100110111110000110111001001010;
		10'd470: 32'b11110111011011010100110111101011;
		10'd471: 32'b00111111001001100110111100110000;
		10'd472: 32'b01111101101111100110110001111001;
		10'd473: 32'b01100011011011010010101111111001;
		10'd474: 32'b01111101100101000111111010100111;
		10'd475: 32'b01010011011100111110111100100100;
		10'd476: 32'b01101110010001110111111001111101;
		10'd477: 32'b01111001010011101110111011110001;
		10'd478: 32'b00111011010101010110111001111101;
		10'd479: 32'b11111010101111001110111010100100;
		10'd480: 32'b11110010111101001011101101110001;
		10'd481: 32'b11111110001001001110111111000111;
		10'd482: 32'b01111100010100111110101111010011;
		10'd483: 32'b11111010011011111110111010111101;
		10'd484: 32'b10100000111111001111101011110110;
		10'd485: 32'b11111000111011101100101011011010;
		10'd486: 32'b00101110011101011110110111001101;
		10'd487: 32'b11111111011110011000111000101101;
		10'd488: 32'b00100110111011011000111101111110;
		10'd489: 32'b11111001011011111011111000001111;
		10'd490: 32'b11011100111011111001111001110111;
		10'd491: 32'b10101101111000111000111101101111;
		10'd492: 32'b10111110111001101000111001110110;
		10'd493: 32'b10101011111111101000101100111101;
		10'd494: 32'b10101100111001011001110010010011;
		10'd495: 32'b00110101101111110011111101111001;
		10'd496: 32'b11111010011100100101001000101110;
		10'd497: 32'b00110111011011110000011100011100;
		10'd498: 32'b01111110111110101101101110111101;
		10'd499: 32'b00010101011011110111101110011101;
		10'd500: 32'b10110110001011001111000001111100;
		10'd501: 32'b01110111111010111000110011001000;
		10'd502: 32'b10111111001110100110101010111100;
		10'd503: 32'b01111111100101111001111010111111;
		10'd504: 32'b01011111101011111011011111111111;
		10'd505: 32'b11010011101001111101110000010011;
		10'd506: 32'b10110011111111111101000110101011;
		10'd507: 32'b11001110100000110100110001010011;
		10'd508: 32'b10111100111111111101111100110011;
		10'd509: 32'b11110110010100011011110000110011;
		10'd510: 32'b11111110001111111110110100101111;
		10'd511: 32'b11101101011101100010011111111111;
		10'd512: 32'b01010101101100110000111011110010;
		10'd513: 32'b01111111110101010010111110101111;
		10'd514: 32'b11111111101111111101101110111110;
		10'd515: 32'b11101111101101011011111111111111;
		10'd516: 32'b01011001101111110010111110110111;
		10'd517: 32'b01111011110100010100111111111111;
		10'd518: 32'b11110111111101110111111110110111;
		10'd519: 32'b11111101101011011010111101011111;
		10'd520: 32'b10111001101111110001111101101100;
		10'd521: 32'b10111100101011100001111011111001;
		10'd522: 32'b11111101101111101101111110111111;
		10'd523: 32'b00011110111010011110101101110101;
		10'd524: 32'b11011110010111000111110111111110;
		10'd525: 32'b11111001101001111110111111111011;
		10'd526: 32'b11111101101111001101101101111101;
		10'd527: 32'b01110011101011000111010000010110;
		10'd528: 32'b11111011011001101001100111111011;
		10'd529: 32'b11110001000001110111111101111110;
		10'd530: 32'b10110011101101010011100110000010;
		10'd531: 32'b11110011100010111011011101110010;
		10'd532: 32'b01111111011001100101101111111010;
		10'd533: 32'b11111101001111110011011011111111;
		10'd534: 32'b11101001001111111001100111110110;
		10'd535: 32'b11101101111011101111111000111110;
		10'd536: 32'b01110111111101101111110010111110;
		10'd537: 32'b11111110111111101011100100100000;
		10'd538: 32'b01100110101011011010111011110111;
		10'd539: 32'b11101001100111001111111110100111;
		10'd540: 32'b11111110011001011110111011111100;
		10'd541: 32'b11111110011001111110111110010011;
		10'd542: 32'b10111110111110011111111111111111;
		10'd543: 32'b01110000111010011100001111010110;
		10'd544: 32'b00011011110101111110101111111101;
		10'd545: 32'b11111011110100011010110111111111;
		10'd546: 32'b00111111110101100001101001110101;
		10'd547: 32'b01111000111111000100110110001110;
		10'd548: 32'b01011111110101011010100101001101;
		10'd549: 32'b00010101111101000111111110011111;
		10'd550: 32'b00110011110001111101111001001111;
		10'd551: 32'b11101011111111111100111101111000;
		10'd552: 32'b11101011111100111111111110100111;
		10'd553: 32'b00101001111110111010110100111100;
		10'd554: 32'b11100011110110001010110111100011;
		10'd555: 32'b11011001101110110101111001111101;
		10'd556: 32'b11101111111111111110101111001111;
		10'd557: 32'b01101011110111101110111101111101;
		10'd558: 32'b11011011011111111110110111101110;
		10'd559: 32'b11111000110111110111100011011100;
		10'd560: 32'b11101010111101100111001011010110;
		10'd561: 32'b01111011111100111001000111111111;
		10'd562: 32'b00101010101111111101101011101101;
		10'd563: 32'b11111001111111111011100111101101;
		10'd564: 32'b01111010101100101110001011111100;
		10'd565: 32'b00001111111000111011100011101111;
		10'd566: 32'b00101100101111111001100011110111;
		10'd567: 32'b10100111111111000010010011110100;
		10'd568: 32'b01111111100011110101111111101101;
		10'd569: 32'b10111111110011111101110111110101;
		10'd570: 32'b01101101011000010001111111010110;
		10'd571: 32'b11110111111111100100001010100100;
		10'd572: 32'b00111011010010011001110111110111;
		10'd573: 32'b00111101111011111111011111001101;
		10'd574: 32'b11111010110111011101111011010101;
	endcase;
	return out;
endfunction
