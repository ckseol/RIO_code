package xorshift_rng_r12_m5_logic;
import Vector::*;
(* noinline *)
function Vector#(64, Bit#(32)) parallel_randint32(Bit#(384) x);
	Vector#(64, Bit#(32)) y = replicate(0);
	y[0]=randint0(x);
	y[1]=randint1(x);
	y[2]=randint2(x);
	y[3]=randint3(x);
	y[4]=randint4(x);
	y[5]=randint5(x);
	y[6]=randint6(x);
	y[7]=randint7(x);
	y[8]=randint8(x);
	y[9]=randint9(x);
	y[10]=randint10(x);
	y[11]=randint11(x);
	y[12]=randint12(x);
	y[13]=randint13(x);
	y[14]=randint14(x);
	y[15]=randint15(x);
	y[16]=randint16(x);
	y[17]=randint17(x);
	y[18]=randint18(x);
	y[19]=randint19(x);
	y[20]=randint20(x);
	y[21]=randint21(x);
	y[22]=randint22(x);
	y[23]=randint23(x);
	y[24]=randint24(x);
	y[25]=randint25(x);
	y[26]=randint26(x);
	y[27]=randint27(x);
	y[28]=randint28(x);
	y[29]=randint29(x);
	y[30]=randint30(x);
	y[31]=randint31(x);
	y[32]=randint32(x);
	y[33]=randint33(x);
	y[34]=randint34(x);
	y[35]=randint35(x);
	y[36]=randint36(x);
	y[37]=randint37(x);
	y[38]=randint38(x);
	y[39]=randint39(x);
	y[40]=randint40(x);
	y[41]=randint41(x);
	y[42]=randint42(x);
	y[43]=randint43(x);
	y[44]=randint44(x);
	y[45]=randint45(x);
	y[46]=randint46(x);
	y[47]=randint47(x);
	y[48]=randint48(x);
	y[49]=randint49(x);
	y[50]=randint50(x);
	y[51]=randint51(x);
	y[52]=randint52(x);
	y[53]=randint53(x);
	y[54]=randint54(x);
	y[55]=randint55(x);
	y[56]=randint56(x);
	y[57]=randint57(x);
	y[58]=randint58(x);
	y[59]=randint59(x);
	y[60]=randint60(x);
	y[61]=randint61(x);
	y[62]=randint62(x);
	y[63]=randint63(x);
	return y;
endfunction

(* noinline *)
function Bit#(32) randint0(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[373]^x[362]^x[159]^x[153];
	y[30]=x[382]^x[372]^x[361]^x[158]^x[152];
	y[29]=x[381]^x[371]^x[360]^x[157]^x[151];
	y[28]=x[380]^x[370]^x[359]^x[156]^x[150];
	y[27]=x[379]^x[369]^x[358]^x[155]^x[149];
	y[26]=x[378]^x[368]^x[357]^x[154]^x[148];
	y[25]=x[377]^x[367]^x[356]^x[153]^x[147];
	y[24]=x[376]^x[366]^x[355]^x[152]^x[146];
	y[23]=x[375]^x[365]^x[354]^x[151]^x[145];
	y[22]=x[374]^x[364]^x[353]^x[150]^x[144];
	y[21]=x[373]^x[363]^x[352]^x[149]^x[143];
	y[20]=x[383]^x[372]^x[148]^x[142];
	y[19]=x[382]^x[371]^x[147]^x[141];
	y[18]=x[381]^x[370]^x[146]^x[140];
	y[17]=x[380]^x[369]^x[145]^x[139];
	y[16]=x[379]^x[368]^x[144]^x[138];
	y[15]=x[378]^x[367]^x[143]^x[137];
	y[14]=x[377]^x[366]^x[142]^x[136];
	y[13]=x[376]^x[365]^x[141]^x[135];
	y[12]=x[375]^x[364]^x[140]^x[134];
	y[11]=x[374]^x[363]^x[139]^x[133];
	y[10]=x[373]^x[362]^x[138]^x[132];
	y[9]=x[372]^x[361]^x[137]^x[131];
	y[8]=x[371]^x[360]^x[136]^x[130];
	y[7]=x[370]^x[359]^x[135]^x[129];
	y[6]=x[369]^x[358]^x[134]^x[128];
	y[5]=x[368]^x[357]^x[133];
	y[4]=x[367]^x[356]^x[132];
	y[3]=x[366]^x[355]^x[131];
	y[2]=x[365]^x[354]^x[130];
	y[1]=x[364]^x[353]^x[129];
	y[0]=x[363]^x[352]^x[128];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint1(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[341]^x[330]^x[127]^x[121];
	y[30]=x[350]^x[340]^x[329]^x[126]^x[120];
	y[29]=x[349]^x[339]^x[328]^x[125]^x[119];
	y[28]=x[348]^x[338]^x[327]^x[124]^x[118];
	y[27]=x[347]^x[337]^x[326]^x[123]^x[117];
	y[26]=x[346]^x[336]^x[325]^x[122]^x[116];
	y[25]=x[345]^x[335]^x[324]^x[121]^x[115];
	y[24]=x[344]^x[334]^x[323]^x[120]^x[114];
	y[23]=x[343]^x[333]^x[322]^x[119]^x[113];
	y[22]=x[342]^x[332]^x[321]^x[118]^x[112];
	y[21]=x[341]^x[331]^x[320]^x[117]^x[111];
	y[20]=x[351]^x[340]^x[116]^x[110];
	y[19]=x[350]^x[339]^x[115]^x[109];
	y[18]=x[349]^x[338]^x[114]^x[108];
	y[17]=x[348]^x[337]^x[113]^x[107];
	y[16]=x[347]^x[336]^x[112]^x[106];
	y[15]=x[346]^x[335]^x[111]^x[105];
	y[14]=x[345]^x[334]^x[110]^x[104];
	y[13]=x[344]^x[333]^x[109]^x[103];
	y[12]=x[343]^x[332]^x[108]^x[102];
	y[11]=x[342]^x[331]^x[107]^x[101];
	y[10]=x[341]^x[330]^x[106]^x[100];
	y[9]=x[340]^x[329]^x[105]^x[99];
	y[8]=x[339]^x[328]^x[104]^x[98];
	y[7]=x[338]^x[327]^x[103]^x[97];
	y[6]=x[337]^x[326]^x[102]^x[96];
	y[5]=x[336]^x[325]^x[101];
	y[4]=x[335]^x[324]^x[100];
	y[3]=x[334]^x[323]^x[99];
	y[2]=x[333]^x[322]^x[98];
	y[1]=x[332]^x[321]^x[97];
	y[0]=x[331]^x[320]^x[96];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint2(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[319]^x[309]^x[298]^x[95]^x[89];
	y[30]=x[318]^x[308]^x[297]^x[94]^x[88];
	y[29]=x[317]^x[307]^x[296]^x[93]^x[87];
	y[28]=x[316]^x[306]^x[295]^x[92]^x[86];
	y[27]=x[315]^x[305]^x[294]^x[91]^x[85];
	y[26]=x[314]^x[304]^x[293]^x[90]^x[84];
	y[25]=x[313]^x[303]^x[292]^x[89]^x[83];
	y[24]=x[312]^x[302]^x[291]^x[88]^x[82];
	y[23]=x[311]^x[301]^x[290]^x[87]^x[81];
	y[22]=x[310]^x[300]^x[289]^x[86]^x[80];
	y[21]=x[309]^x[299]^x[288]^x[85]^x[79];
	y[20]=x[319]^x[308]^x[84]^x[78];
	y[19]=x[318]^x[307]^x[83]^x[77];
	y[18]=x[317]^x[306]^x[82]^x[76];
	y[17]=x[316]^x[305]^x[81]^x[75];
	y[16]=x[315]^x[304]^x[80]^x[74];
	y[15]=x[314]^x[303]^x[79]^x[73];
	y[14]=x[313]^x[302]^x[78]^x[72];
	y[13]=x[312]^x[301]^x[77]^x[71];
	y[12]=x[311]^x[300]^x[76]^x[70];
	y[11]=x[310]^x[299]^x[75]^x[69];
	y[10]=x[309]^x[298]^x[74]^x[68];
	y[9]=x[308]^x[297]^x[73]^x[67];
	y[8]=x[307]^x[296]^x[72]^x[66];
	y[7]=x[306]^x[295]^x[71]^x[65];
	y[6]=x[305]^x[294]^x[70]^x[64];
	y[5]=x[304]^x[293]^x[69];
	y[4]=x[303]^x[292]^x[68];
	y[3]=x[302]^x[291]^x[67];
	y[2]=x[301]^x[290]^x[66];
	y[1]=x[300]^x[289]^x[65];
	y[0]=x[299]^x[288]^x[64];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint3(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[287]^x[277]^x[266]^x[63]^x[57];
	y[30]=x[286]^x[276]^x[265]^x[62]^x[56];
	y[29]=x[285]^x[275]^x[264]^x[61]^x[55];
	y[28]=x[284]^x[274]^x[263]^x[60]^x[54];
	y[27]=x[283]^x[273]^x[262]^x[59]^x[53];
	y[26]=x[282]^x[272]^x[261]^x[58]^x[52];
	y[25]=x[281]^x[271]^x[260]^x[57]^x[51];
	y[24]=x[280]^x[270]^x[259]^x[56]^x[50];
	y[23]=x[279]^x[269]^x[258]^x[55]^x[49];
	y[22]=x[278]^x[268]^x[257]^x[54]^x[48];
	y[21]=x[277]^x[267]^x[256]^x[53]^x[47];
	y[20]=x[287]^x[276]^x[52]^x[46];
	y[19]=x[286]^x[275]^x[51]^x[45];
	y[18]=x[285]^x[274]^x[50]^x[44];
	y[17]=x[284]^x[273]^x[49]^x[43];
	y[16]=x[283]^x[272]^x[48]^x[42];
	y[15]=x[282]^x[271]^x[47]^x[41];
	y[14]=x[281]^x[270]^x[46]^x[40];
	y[13]=x[280]^x[269]^x[45]^x[39];
	y[12]=x[279]^x[268]^x[44]^x[38];
	y[11]=x[278]^x[267]^x[43]^x[37];
	y[10]=x[277]^x[266]^x[42]^x[36];
	y[9]=x[276]^x[265]^x[41]^x[35];
	y[8]=x[275]^x[264]^x[40]^x[34];
	y[7]=x[274]^x[263]^x[39]^x[33];
	y[6]=x[273]^x[262]^x[38]^x[32];
	y[5]=x[272]^x[261]^x[37];
	y[4]=x[271]^x[260]^x[36];
	y[3]=x[270]^x[259]^x[35];
	y[2]=x[269]^x[258]^x[34];
	y[1]=x[268]^x[257]^x[33];
	y[0]=x[267]^x[256]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint4(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[255]^x[245]^x[234]^x[31]^x[25];
	y[30]=x[254]^x[244]^x[233]^x[30]^x[24];
	y[29]=x[253]^x[243]^x[232]^x[29]^x[23];
	y[28]=x[252]^x[242]^x[231]^x[28]^x[22];
	y[27]=x[251]^x[241]^x[230]^x[27]^x[21];
	y[26]=x[250]^x[240]^x[229]^x[26]^x[20];
	y[25]=x[249]^x[239]^x[228]^x[25]^x[19];
	y[24]=x[248]^x[238]^x[227]^x[24]^x[18];
	y[23]=x[247]^x[237]^x[226]^x[23]^x[17];
	y[22]=x[246]^x[236]^x[225]^x[22]^x[16];
	y[21]=x[245]^x[235]^x[224]^x[21]^x[15];
	y[20]=x[255]^x[244]^x[20]^x[14];
	y[19]=x[254]^x[243]^x[19]^x[13];
	y[18]=x[253]^x[242]^x[18]^x[12];
	y[17]=x[252]^x[241]^x[17]^x[11];
	y[16]=x[251]^x[240]^x[16]^x[10];
	y[15]=x[250]^x[239]^x[15]^x[9];
	y[14]=x[249]^x[238]^x[14]^x[8];
	y[13]=x[248]^x[237]^x[13]^x[7];
	y[12]=x[247]^x[236]^x[12]^x[6];
	y[11]=x[246]^x[235]^x[11]^x[5];
	y[10]=x[245]^x[234]^x[10]^x[4];
	y[9]=x[244]^x[233]^x[9]^x[3];
	y[8]=x[243]^x[232]^x[8]^x[2];
	y[7]=x[242]^x[231]^x[7]^x[1];
	y[6]=x[241]^x[230]^x[6]^x[0];
	y[5]=x[240]^x[229]^x[5];
	y[4]=x[239]^x[228]^x[4];
	y[3]=x[238]^x[227]^x[3];
	y[2]=x[237]^x[226]^x[2];
	y[1]=x[236]^x[225]^x[1];
	y[0]=x[235]^x[224]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint5(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[377]^x[373]^x[367]^x[362]^x[356]^x[223]^x[213]^x[202]^x[159]^x[147];
	y[30]=x[382]^x[376]^x[372]^x[366]^x[361]^x[355]^x[222]^x[212]^x[201]^x[158]^x[146];
	y[29]=x[381]^x[375]^x[371]^x[365]^x[360]^x[354]^x[221]^x[211]^x[200]^x[157]^x[145];
	y[28]=x[380]^x[374]^x[370]^x[364]^x[359]^x[353]^x[220]^x[210]^x[199]^x[156]^x[144];
	y[27]=x[379]^x[373]^x[369]^x[363]^x[358]^x[352]^x[219]^x[209]^x[198]^x[155]^x[143];
	y[26]=x[383]^x[378]^x[372]^x[368]^x[357]^x[218]^x[208]^x[197]^x[154]^x[142];
	y[25]=x[382]^x[377]^x[371]^x[367]^x[356]^x[217]^x[207]^x[196]^x[153]^x[141];
	y[24]=x[381]^x[376]^x[370]^x[366]^x[355]^x[216]^x[206]^x[195]^x[152]^x[140];
	y[23]=x[380]^x[375]^x[369]^x[365]^x[354]^x[215]^x[205]^x[194]^x[151]^x[139];
	y[22]=x[379]^x[374]^x[368]^x[364]^x[353]^x[214]^x[204]^x[193]^x[150]^x[138];
	y[21]=x[378]^x[373]^x[367]^x[363]^x[352]^x[213]^x[203]^x[192]^x[149]^x[137];
	y[20]=x[383]^x[377]^x[372]^x[366]^x[223]^x[212]^x[148]^x[136];
	y[19]=x[382]^x[376]^x[371]^x[365]^x[222]^x[211]^x[147]^x[135];
	y[18]=x[381]^x[375]^x[370]^x[364]^x[221]^x[210]^x[146]^x[134];
	y[17]=x[380]^x[374]^x[369]^x[363]^x[220]^x[209]^x[145]^x[133];
	y[16]=x[379]^x[373]^x[368]^x[362]^x[219]^x[208]^x[144]^x[132];
	y[15]=x[378]^x[372]^x[367]^x[361]^x[218]^x[207]^x[143]^x[131];
	y[14]=x[377]^x[371]^x[366]^x[360]^x[217]^x[206]^x[142]^x[130];
	y[13]=x[376]^x[370]^x[365]^x[359]^x[216]^x[205]^x[141]^x[129];
	y[12]=x[375]^x[369]^x[364]^x[358]^x[215]^x[204]^x[140]^x[128];
	y[11]=x[374]^x[368]^x[363]^x[357]^x[214]^x[203]^x[139];
	y[10]=x[373]^x[367]^x[362]^x[356]^x[213]^x[202]^x[138];
	y[9]=x[372]^x[366]^x[361]^x[355]^x[212]^x[201]^x[137];
	y[8]=x[371]^x[365]^x[360]^x[354]^x[211]^x[200]^x[136];
	y[7]=x[370]^x[364]^x[359]^x[353]^x[210]^x[199]^x[135];
	y[6]=x[369]^x[363]^x[358]^x[352]^x[209]^x[198]^x[134];
	y[5]=x[368]^x[357]^x[208]^x[197]^x[133];
	y[4]=x[367]^x[356]^x[207]^x[196]^x[132];
	y[3]=x[366]^x[355]^x[206]^x[195]^x[131];
	y[2]=x[365]^x[354]^x[205]^x[194]^x[130];
	y[1]=x[364]^x[353]^x[204]^x[193]^x[129];
	y[0]=x[363]^x[352]^x[203]^x[192]^x[128];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint6(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[345]^x[341]^x[335]^x[330]^x[324]^x[191]^x[181]^x[170]^x[127]^x[115];
	y[30]=x[350]^x[344]^x[340]^x[334]^x[329]^x[323]^x[190]^x[180]^x[169]^x[126]^x[114];
	y[29]=x[349]^x[343]^x[339]^x[333]^x[328]^x[322]^x[189]^x[179]^x[168]^x[125]^x[113];
	y[28]=x[348]^x[342]^x[338]^x[332]^x[327]^x[321]^x[188]^x[178]^x[167]^x[124]^x[112];
	y[27]=x[347]^x[341]^x[337]^x[331]^x[326]^x[320]^x[187]^x[177]^x[166]^x[123]^x[111];
	y[26]=x[351]^x[346]^x[340]^x[336]^x[325]^x[186]^x[176]^x[165]^x[122]^x[110];
	y[25]=x[350]^x[345]^x[339]^x[335]^x[324]^x[185]^x[175]^x[164]^x[121]^x[109];
	y[24]=x[349]^x[344]^x[338]^x[334]^x[323]^x[184]^x[174]^x[163]^x[120]^x[108];
	y[23]=x[348]^x[343]^x[337]^x[333]^x[322]^x[183]^x[173]^x[162]^x[119]^x[107];
	y[22]=x[347]^x[342]^x[336]^x[332]^x[321]^x[182]^x[172]^x[161]^x[118]^x[106];
	y[21]=x[346]^x[341]^x[335]^x[331]^x[320]^x[181]^x[171]^x[160]^x[117]^x[105];
	y[20]=x[351]^x[345]^x[340]^x[334]^x[191]^x[180]^x[116]^x[104];
	y[19]=x[350]^x[344]^x[339]^x[333]^x[190]^x[179]^x[115]^x[103];
	y[18]=x[349]^x[343]^x[338]^x[332]^x[189]^x[178]^x[114]^x[102];
	y[17]=x[348]^x[342]^x[337]^x[331]^x[188]^x[177]^x[113]^x[101];
	y[16]=x[347]^x[341]^x[336]^x[330]^x[187]^x[176]^x[112]^x[100];
	y[15]=x[346]^x[340]^x[335]^x[329]^x[186]^x[175]^x[111]^x[99];
	y[14]=x[345]^x[339]^x[334]^x[328]^x[185]^x[174]^x[110]^x[98];
	y[13]=x[344]^x[338]^x[333]^x[327]^x[184]^x[173]^x[109]^x[97];
	y[12]=x[343]^x[337]^x[332]^x[326]^x[183]^x[172]^x[108]^x[96];
	y[11]=x[342]^x[336]^x[331]^x[325]^x[182]^x[171]^x[107];
	y[10]=x[341]^x[335]^x[330]^x[324]^x[181]^x[170]^x[106];
	y[9]=x[340]^x[334]^x[329]^x[323]^x[180]^x[169]^x[105];
	y[8]=x[339]^x[333]^x[328]^x[322]^x[179]^x[168]^x[104];
	y[7]=x[338]^x[332]^x[327]^x[321]^x[178]^x[167]^x[103];
	y[6]=x[337]^x[331]^x[326]^x[320]^x[177]^x[166]^x[102];
	y[5]=x[336]^x[325]^x[176]^x[165]^x[101];
	y[4]=x[335]^x[324]^x[175]^x[164]^x[100];
	y[3]=x[334]^x[323]^x[174]^x[163]^x[99];
	y[2]=x[333]^x[322]^x[173]^x[162]^x[98];
	y[1]=x[332]^x[321]^x[172]^x[161]^x[97];
	y[0]=x[331]^x[320]^x[171]^x[160]^x[96];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint7(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[319]^x[313]^x[309]^x[303]^x[298]^x[292]^x[159]^x[149]^x[138]^x[95]^x[83];
	y[30]=x[318]^x[312]^x[308]^x[302]^x[297]^x[291]^x[158]^x[148]^x[137]^x[94]^x[82];
	y[29]=x[317]^x[311]^x[307]^x[301]^x[296]^x[290]^x[157]^x[147]^x[136]^x[93]^x[81];
	y[28]=x[316]^x[310]^x[306]^x[300]^x[295]^x[289]^x[156]^x[146]^x[135]^x[92]^x[80];
	y[27]=x[315]^x[309]^x[305]^x[299]^x[294]^x[288]^x[155]^x[145]^x[134]^x[91]^x[79];
	y[26]=x[319]^x[314]^x[308]^x[304]^x[293]^x[154]^x[144]^x[133]^x[90]^x[78];
	y[25]=x[318]^x[313]^x[307]^x[303]^x[292]^x[153]^x[143]^x[132]^x[89]^x[77];
	y[24]=x[317]^x[312]^x[306]^x[302]^x[291]^x[152]^x[142]^x[131]^x[88]^x[76];
	y[23]=x[316]^x[311]^x[305]^x[301]^x[290]^x[151]^x[141]^x[130]^x[87]^x[75];
	y[22]=x[315]^x[310]^x[304]^x[300]^x[289]^x[150]^x[140]^x[129]^x[86]^x[74];
	y[21]=x[314]^x[309]^x[303]^x[299]^x[288]^x[149]^x[139]^x[128]^x[85]^x[73];
	y[20]=x[319]^x[313]^x[308]^x[302]^x[159]^x[148]^x[84]^x[72];
	y[19]=x[318]^x[312]^x[307]^x[301]^x[158]^x[147]^x[83]^x[71];
	y[18]=x[317]^x[311]^x[306]^x[300]^x[157]^x[146]^x[82]^x[70];
	y[17]=x[316]^x[310]^x[305]^x[299]^x[156]^x[145]^x[81]^x[69];
	y[16]=x[315]^x[309]^x[304]^x[298]^x[155]^x[144]^x[80]^x[68];
	y[15]=x[314]^x[308]^x[303]^x[297]^x[154]^x[143]^x[79]^x[67];
	y[14]=x[313]^x[307]^x[302]^x[296]^x[153]^x[142]^x[78]^x[66];
	y[13]=x[312]^x[306]^x[301]^x[295]^x[152]^x[141]^x[77]^x[65];
	y[12]=x[311]^x[305]^x[300]^x[294]^x[151]^x[140]^x[76]^x[64];
	y[11]=x[310]^x[304]^x[299]^x[293]^x[150]^x[139]^x[75];
	y[10]=x[309]^x[303]^x[298]^x[292]^x[149]^x[138]^x[74];
	y[9]=x[308]^x[302]^x[297]^x[291]^x[148]^x[137]^x[73];
	y[8]=x[307]^x[301]^x[296]^x[290]^x[147]^x[136]^x[72];
	y[7]=x[306]^x[300]^x[295]^x[289]^x[146]^x[135]^x[71];
	y[6]=x[305]^x[299]^x[294]^x[288]^x[145]^x[134]^x[70];
	y[5]=x[304]^x[293]^x[144]^x[133]^x[69];
	y[4]=x[303]^x[292]^x[143]^x[132]^x[68];
	y[3]=x[302]^x[291]^x[142]^x[131]^x[67];
	y[2]=x[301]^x[290]^x[141]^x[130]^x[66];
	y[1]=x[300]^x[289]^x[140]^x[129]^x[65];
	y[0]=x[299]^x[288]^x[139]^x[128]^x[64];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint8(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[287]^x[281]^x[277]^x[271]^x[266]^x[260]^x[127]^x[117]^x[106]^x[63]^x[51];
	y[30]=x[286]^x[280]^x[276]^x[270]^x[265]^x[259]^x[126]^x[116]^x[105]^x[62]^x[50];
	y[29]=x[285]^x[279]^x[275]^x[269]^x[264]^x[258]^x[125]^x[115]^x[104]^x[61]^x[49];
	y[28]=x[284]^x[278]^x[274]^x[268]^x[263]^x[257]^x[124]^x[114]^x[103]^x[60]^x[48];
	y[27]=x[283]^x[277]^x[273]^x[267]^x[262]^x[256]^x[123]^x[113]^x[102]^x[59]^x[47];
	y[26]=x[287]^x[282]^x[276]^x[272]^x[261]^x[122]^x[112]^x[101]^x[58]^x[46];
	y[25]=x[286]^x[281]^x[275]^x[271]^x[260]^x[121]^x[111]^x[100]^x[57]^x[45];
	y[24]=x[285]^x[280]^x[274]^x[270]^x[259]^x[120]^x[110]^x[99]^x[56]^x[44];
	y[23]=x[284]^x[279]^x[273]^x[269]^x[258]^x[119]^x[109]^x[98]^x[55]^x[43];
	y[22]=x[283]^x[278]^x[272]^x[268]^x[257]^x[118]^x[108]^x[97]^x[54]^x[42];
	y[21]=x[282]^x[277]^x[271]^x[267]^x[256]^x[117]^x[107]^x[96]^x[53]^x[41];
	y[20]=x[287]^x[281]^x[276]^x[270]^x[127]^x[116]^x[52]^x[40];
	y[19]=x[286]^x[280]^x[275]^x[269]^x[126]^x[115]^x[51]^x[39];
	y[18]=x[285]^x[279]^x[274]^x[268]^x[125]^x[114]^x[50]^x[38];
	y[17]=x[284]^x[278]^x[273]^x[267]^x[124]^x[113]^x[49]^x[37];
	y[16]=x[283]^x[277]^x[272]^x[266]^x[123]^x[112]^x[48]^x[36];
	y[15]=x[282]^x[276]^x[271]^x[265]^x[122]^x[111]^x[47]^x[35];
	y[14]=x[281]^x[275]^x[270]^x[264]^x[121]^x[110]^x[46]^x[34];
	y[13]=x[280]^x[274]^x[269]^x[263]^x[120]^x[109]^x[45]^x[33];
	y[12]=x[279]^x[273]^x[268]^x[262]^x[119]^x[108]^x[44]^x[32];
	y[11]=x[278]^x[272]^x[267]^x[261]^x[118]^x[107]^x[43];
	y[10]=x[277]^x[271]^x[266]^x[260]^x[117]^x[106]^x[42];
	y[9]=x[276]^x[270]^x[265]^x[259]^x[116]^x[105]^x[41];
	y[8]=x[275]^x[269]^x[264]^x[258]^x[115]^x[104]^x[40];
	y[7]=x[274]^x[268]^x[263]^x[257]^x[114]^x[103]^x[39];
	y[6]=x[273]^x[267]^x[262]^x[256]^x[113]^x[102]^x[38];
	y[5]=x[272]^x[261]^x[112]^x[101]^x[37];
	y[4]=x[271]^x[260]^x[111]^x[100]^x[36];
	y[3]=x[270]^x[259]^x[110]^x[99]^x[35];
	y[2]=x[269]^x[258]^x[109]^x[98]^x[34];
	y[1]=x[268]^x[257]^x[108]^x[97]^x[33];
	y[0]=x[267]^x[256]^x[107]^x[96]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint9(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[255]^x[249]^x[245]^x[239]^x[234]^x[228]^x[95]^x[85]^x[74]^x[31]^x[19];
	y[30]=x[254]^x[248]^x[244]^x[238]^x[233]^x[227]^x[94]^x[84]^x[73]^x[30]^x[18];
	y[29]=x[253]^x[247]^x[243]^x[237]^x[232]^x[226]^x[93]^x[83]^x[72]^x[29]^x[17];
	y[28]=x[252]^x[246]^x[242]^x[236]^x[231]^x[225]^x[92]^x[82]^x[71]^x[28]^x[16];
	y[27]=x[251]^x[245]^x[241]^x[235]^x[230]^x[224]^x[91]^x[81]^x[70]^x[27]^x[15];
	y[26]=x[255]^x[250]^x[244]^x[240]^x[229]^x[90]^x[80]^x[69]^x[26]^x[14];
	y[25]=x[254]^x[249]^x[243]^x[239]^x[228]^x[89]^x[79]^x[68]^x[25]^x[13];
	y[24]=x[253]^x[248]^x[242]^x[238]^x[227]^x[88]^x[78]^x[67]^x[24]^x[12];
	y[23]=x[252]^x[247]^x[241]^x[237]^x[226]^x[87]^x[77]^x[66]^x[23]^x[11];
	y[22]=x[251]^x[246]^x[240]^x[236]^x[225]^x[86]^x[76]^x[65]^x[22]^x[10];
	y[21]=x[250]^x[245]^x[239]^x[235]^x[224]^x[85]^x[75]^x[64]^x[21]^x[9];
	y[20]=x[255]^x[249]^x[244]^x[238]^x[95]^x[84]^x[20]^x[8];
	y[19]=x[254]^x[248]^x[243]^x[237]^x[94]^x[83]^x[19]^x[7];
	y[18]=x[253]^x[247]^x[242]^x[236]^x[93]^x[82]^x[18]^x[6];
	y[17]=x[252]^x[246]^x[241]^x[235]^x[92]^x[81]^x[17]^x[5];
	y[16]=x[251]^x[245]^x[240]^x[234]^x[91]^x[80]^x[16]^x[4];
	y[15]=x[250]^x[244]^x[239]^x[233]^x[90]^x[79]^x[15]^x[3];
	y[14]=x[249]^x[243]^x[238]^x[232]^x[89]^x[78]^x[14]^x[2];
	y[13]=x[248]^x[242]^x[237]^x[231]^x[88]^x[77]^x[13]^x[1];
	y[12]=x[247]^x[241]^x[236]^x[230]^x[87]^x[76]^x[12]^x[0];
	y[11]=x[246]^x[240]^x[235]^x[229]^x[86]^x[75]^x[11];
	y[10]=x[245]^x[239]^x[234]^x[228]^x[85]^x[74]^x[10];
	y[9]=x[244]^x[238]^x[233]^x[227]^x[84]^x[73]^x[9];
	y[8]=x[243]^x[237]^x[232]^x[226]^x[83]^x[72]^x[8];
	y[7]=x[242]^x[236]^x[231]^x[225]^x[82]^x[71]^x[7];
	y[6]=x[241]^x[235]^x[230]^x[224]^x[81]^x[70]^x[6];
	y[5]=x[240]^x[229]^x[80]^x[69]^x[5];
	y[4]=x[239]^x[228]^x[79]^x[68]^x[4];
	y[3]=x[238]^x[227]^x[78]^x[67]^x[3];
	y[2]=x[237]^x[226]^x[77]^x[66]^x[2];
	y[1]=x[236]^x[225]^x[76]^x[65]^x[1];
	y[0]=x[235]^x[224]^x[75]^x[64]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint10(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[373]^x[371]^x[362]^x[223]^x[217]^x[213]^x[207]^x[202]^x[196]^x[159]^x[153]^x[147]^x[141]^x[63]^x[53]^x[42];
	y[30]=x[382]^x[381]^x[372]^x[370]^x[361]^x[222]^x[216]^x[212]^x[206]^x[201]^x[195]^x[158]^x[152]^x[146]^x[140]^x[62]^x[52]^x[41];
	y[29]=x[381]^x[380]^x[371]^x[369]^x[360]^x[221]^x[215]^x[211]^x[205]^x[200]^x[194]^x[157]^x[151]^x[145]^x[139]^x[61]^x[51]^x[40];
	y[28]=x[380]^x[379]^x[370]^x[368]^x[359]^x[220]^x[214]^x[210]^x[204]^x[199]^x[193]^x[156]^x[150]^x[144]^x[138]^x[60]^x[50]^x[39];
	y[27]=x[379]^x[378]^x[369]^x[367]^x[358]^x[219]^x[213]^x[209]^x[203]^x[198]^x[192]^x[155]^x[149]^x[143]^x[137]^x[59]^x[49]^x[38];
	y[26]=x[378]^x[377]^x[368]^x[366]^x[357]^x[223]^x[218]^x[212]^x[208]^x[197]^x[154]^x[148]^x[142]^x[136]^x[58]^x[48]^x[37];
	y[25]=x[377]^x[376]^x[367]^x[365]^x[356]^x[222]^x[217]^x[211]^x[207]^x[196]^x[153]^x[147]^x[141]^x[135]^x[57]^x[47]^x[36];
	y[24]=x[376]^x[375]^x[366]^x[364]^x[355]^x[221]^x[216]^x[210]^x[206]^x[195]^x[152]^x[146]^x[140]^x[134]^x[56]^x[46]^x[35];
	y[23]=x[375]^x[374]^x[365]^x[363]^x[354]^x[220]^x[215]^x[209]^x[205]^x[194]^x[151]^x[145]^x[139]^x[133]^x[55]^x[45]^x[34];
	y[22]=x[374]^x[373]^x[364]^x[362]^x[353]^x[219]^x[214]^x[208]^x[204]^x[193]^x[150]^x[144]^x[138]^x[132]^x[54]^x[44]^x[33];
	y[21]=x[373]^x[372]^x[363]^x[361]^x[352]^x[218]^x[213]^x[207]^x[203]^x[192]^x[149]^x[143]^x[137]^x[131]^x[53]^x[43]^x[32];
	y[20]=x[383]^x[372]^x[371]^x[360]^x[223]^x[217]^x[212]^x[206]^x[148]^x[142]^x[136]^x[130]^x[63]^x[52];
	y[19]=x[382]^x[371]^x[370]^x[359]^x[222]^x[216]^x[211]^x[205]^x[147]^x[141]^x[135]^x[129]^x[62]^x[51];
	y[18]=x[381]^x[370]^x[369]^x[358]^x[221]^x[215]^x[210]^x[204]^x[146]^x[140]^x[134]^x[128]^x[61]^x[50];
	y[17]=x[380]^x[369]^x[368]^x[357]^x[220]^x[214]^x[209]^x[203]^x[145]^x[139]^x[133]^x[60]^x[49];
	y[16]=x[379]^x[368]^x[367]^x[356]^x[219]^x[213]^x[208]^x[202]^x[144]^x[138]^x[132]^x[59]^x[48];
	y[15]=x[378]^x[367]^x[366]^x[355]^x[218]^x[212]^x[207]^x[201]^x[143]^x[137]^x[131]^x[58]^x[47];
	y[14]=x[377]^x[366]^x[365]^x[354]^x[217]^x[211]^x[206]^x[200]^x[142]^x[136]^x[130]^x[57]^x[46];
	y[13]=x[376]^x[365]^x[364]^x[353]^x[216]^x[210]^x[205]^x[199]^x[141]^x[135]^x[129]^x[56]^x[45];
	y[12]=x[375]^x[364]^x[363]^x[352]^x[215]^x[209]^x[204]^x[198]^x[140]^x[134]^x[128]^x[55]^x[44];
	y[11]=x[374]^x[363]^x[214]^x[208]^x[203]^x[197]^x[139]^x[133]^x[54]^x[43];
	y[10]=x[373]^x[362]^x[213]^x[207]^x[202]^x[196]^x[138]^x[132]^x[53]^x[42];
	y[9]=x[372]^x[361]^x[212]^x[206]^x[201]^x[195]^x[137]^x[131]^x[52]^x[41];
	y[8]=x[371]^x[360]^x[211]^x[205]^x[200]^x[194]^x[136]^x[130]^x[51]^x[40];
	y[7]=x[370]^x[359]^x[210]^x[204]^x[199]^x[193]^x[135]^x[129]^x[50]^x[39];
	y[6]=x[369]^x[358]^x[209]^x[203]^x[198]^x[192]^x[134]^x[128]^x[49]^x[38];
	y[5]=x[368]^x[357]^x[208]^x[197]^x[133]^x[48]^x[37];
	y[4]=x[367]^x[356]^x[207]^x[196]^x[132]^x[47]^x[36];
	y[3]=x[366]^x[355]^x[206]^x[195]^x[131]^x[46]^x[35];
	y[2]=x[365]^x[354]^x[205]^x[194]^x[130]^x[45]^x[34];
	y[1]=x[364]^x[353]^x[204]^x[193]^x[129]^x[44]^x[33];
	y[0]=x[363]^x[352]^x[203]^x[192]^x[128]^x[43]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint11(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[350]^x[341]^x[339]^x[330]^x[191]^x[185]^x[181]^x[175]^x[170]^x[164]^x[127]^x[121]^x[115]^x[109]^x[31]^x[21]^x[10];
	y[30]=x[350]^x[349]^x[340]^x[338]^x[329]^x[190]^x[184]^x[180]^x[174]^x[169]^x[163]^x[126]^x[120]^x[114]^x[108]^x[30]^x[20]^x[9];
	y[29]=x[349]^x[348]^x[339]^x[337]^x[328]^x[189]^x[183]^x[179]^x[173]^x[168]^x[162]^x[125]^x[119]^x[113]^x[107]^x[29]^x[19]^x[8];
	y[28]=x[348]^x[347]^x[338]^x[336]^x[327]^x[188]^x[182]^x[178]^x[172]^x[167]^x[161]^x[124]^x[118]^x[112]^x[106]^x[28]^x[18]^x[7];
	y[27]=x[347]^x[346]^x[337]^x[335]^x[326]^x[187]^x[181]^x[177]^x[171]^x[166]^x[160]^x[123]^x[117]^x[111]^x[105]^x[27]^x[17]^x[6];
	y[26]=x[346]^x[345]^x[336]^x[334]^x[325]^x[191]^x[186]^x[180]^x[176]^x[165]^x[122]^x[116]^x[110]^x[104]^x[26]^x[16]^x[5];
	y[25]=x[345]^x[344]^x[335]^x[333]^x[324]^x[190]^x[185]^x[179]^x[175]^x[164]^x[121]^x[115]^x[109]^x[103]^x[25]^x[15]^x[4];
	y[24]=x[344]^x[343]^x[334]^x[332]^x[323]^x[189]^x[184]^x[178]^x[174]^x[163]^x[120]^x[114]^x[108]^x[102]^x[24]^x[14]^x[3];
	y[23]=x[343]^x[342]^x[333]^x[331]^x[322]^x[188]^x[183]^x[177]^x[173]^x[162]^x[119]^x[113]^x[107]^x[101]^x[23]^x[13]^x[2];
	y[22]=x[342]^x[341]^x[332]^x[330]^x[321]^x[187]^x[182]^x[176]^x[172]^x[161]^x[118]^x[112]^x[106]^x[100]^x[22]^x[12]^x[1];
	y[21]=x[341]^x[340]^x[331]^x[329]^x[320]^x[186]^x[181]^x[175]^x[171]^x[160]^x[117]^x[111]^x[105]^x[99]^x[21]^x[11]^x[0];
	y[20]=x[351]^x[340]^x[339]^x[328]^x[191]^x[185]^x[180]^x[174]^x[116]^x[110]^x[104]^x[98]^x[31]^x[20];
	y[19]=x[350]^x[339]^x[338]^x[327]^x[190]^x[184]^x[179]^x[173]^x[115]^x[109]^x[103]^x[97]^x[30]^x[19];
	y[18]=x[349]^x[338]^x[337]^x[326]^x[189]^x[183]^x[178]^x[172]^x[114]^x[108]^x[102]^x[96]^x[29]^x[18];
	y[17]=x[348]^x[337]^x[336]^x[325]^x[188]^x[182]^x[177]^x[171]^x[113]^x[107]^x[101]^x[28]^x[17];
	y[16]=x[347]^x[336]^x[335]^x[324]^x[187]^x[181]^x[176]^x[170]^x[112]^x[106]^x[100]^x[27]^x[16];
	y[15]=x[346]^x[335]^x[334]^x[323]^x[186]^x[180]^x[175]^x[169]^x[111]^x[105]^x[99]^x[26]^x[15];
	y[14]=x[345]^x[334]^x[333]^x[322]^x[185]^x[179]^x[174]^x[168]^x[110]^x[104]^x[98]^x[25]^x[14];
	y[13]=x[344]^x[333]^x[332]^x[321]^x[184]^x[178]^x[173]^x[167]^x[109]^x[103]^x[97]^x[24]^x[13];
	y[12]=x[343]^x[332]^x[331]^x[320]^x[183]^x[177]^x[172]^x[166]^x[108]^x[102]^x[96]^x[23]^x[12];
	y[11]=x[342]^x[331]^x[182]^x[176]^x[171]^x[165]^x[107]^x[101]^x[22]^x[11];
	y[10]=x[341]^x[330]^x[181]^x[175]^x[170]^x[164]^x[106]^x[100]^x[21]^x[10];
	y[9]=x[340]^x[329]^x[180]^x[174]^x[169]^x[163]^x[105]^x[99]^x[20]^x[9];
	y[8]=x[339]^x[328]^x[179]^x[173]^x[168]^x[162]^x[104]^x[98]^x[19]^x[8];
	y[7]=x[338]^x[327]^x[178]^x[172]^x[167]^x[161]^x[103]^x[97]^x[18]^x[7];
	y[6]=x[337]^x[326]^x[177]^x[171]^x[166]^x[160]^x[102]^x[96]^x[17]^x[6];
	y[5]=x[336]^x[325]^x[176]^x[165]^x[101]^x[16]^x[5];
	y[4]=x[335]^x[324]^x[175]^x[164]^x[100]^x[15]^x[4];
	y[3]=x[334]^x[323]^x[174]^x[163]^x[99]^x[14]^x[3];
	y[2]=x[333]^x[322]^x[173]^x[162]^x[98]^x[13]^x[2];
	y[1]=x[332]^x[321]^x[172]^x[161]^x[97]^x[12]^x[1];
	y[0]=x[331]^x[320]^x[171]^x[160]^x[96]^x[11]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint12(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[373]^x[363]^x[352]^x[319]^x[318]^x[309]^x[307]^x[298]^x[95]^x[89]^x[83]^x[77];
	y[30]=x[383]^x[382]^x[372]^x[318]^x[317]^x[308]^x[306]^x[297]^x[94]^x[88]^x[82]^x[76];
	y[29]=x[382]^x[381]^x[371]^x[317]^x[316]^x[307]^x[305]^x[296]^x[93]^x[87]^x[81]^x[75];
	y[28]=x[381]^x[380]^x[370]^x[316]^x[315]^x[306]^x[304]^x[295]^x[92]^x[86]^x[80]^x[74];
	y[27]=x[380]^x[379]^x[369]^x[315]^x[314]^x[305]^x[303]^x[294]^x[91]^x[85]^x[79]^x[73];
	y[26]=x[379]^x[378]^x[368]^x[314]^x[313]^x[304]^x[302]^x[293]^x[159]^x[138]^x[90]^x[84]^x[78]^x[72];
	y[25]=x[378]^x[377]^x[367]^x[313]^x[312]^x[303]^x[301]^x[292]^x[158]^x[137]^x[89]^x[83]^x[77]^x[71];
	y[24]=x[377]^x[376]^x[366]^x[312]^x[311]^x[302]^x[300]^x[291]^x[157]^x[136]^x[88]^x[82]^x[76]^x[70];
	y[23]=x[376]^x[375]^x[365]^x[311]^x[310]^x[301]^x[299]^x[290]^x[156]^x[135]^x[87]^x[81]^x[75]^x[69];
	y[22]=x[375]^x[374]^x[364]^x[310]^x[309]^x[300]^x[298]^x[289]^x[155]^x[134]^x[86]^x[80]^x[74]^x[68];
	y[21]=x[374]^x[373]^x[363]^x[309]^x[308]^x[299]^x[297]^x[288]^x[154]^x[133]^x[85]^x[79]^x[73]^x[67];
	y[20]=x[373]^x[372]^x[362]^x[319]^x[308]^x[307]^x[296]^x[84]^x[78]^x[72]^x[66];
	y[19]=x[372]^x[371]^x[361]^x[318]^x[307]^x[306]^x[295]^x[83]^x[77]^x[71]^x[65];
	y[18]=x[371]^x[370]^x[360]^x[317]^x[306]^x[305]^x[294]^x[82]^x[76]^x[70]^x[64];
	y[17]=x[370]^x[369]^x[359]^x[316]^x[305]^x[304]^x[293]^x[81]^x[75]^x[69];
	y[16]=x[369]^x[368]^x[358]^x[315]^x[304]^x[303]^x[292]^x[80]^x[74]^x[68];
	y[15]=x[368]^x[367]^x[357]^x[314]^x[303]^x[302]^x[291]^x[79]^x[73]^x[67];
	y[14]=x[367]^x[366]^x[356]^x[313]^x[302]^x[301]^x[290]^x[78]^x[72]^x[66];
	y[13]=x[366]^x[365]^x[355]^x[312]^x[301]^x[300]^x[289]^x[77]^x[71]^x[65];
	y[12]=x[365]^x[364]^x[354]^x[311]^x[300]^x[299]^x[288]^x[76]^x[70]^x[64];
	y[11]=x[364]^x[363]^x[353]^x[310]^x[299]^x[75]^x[69];
	y[10]=x[363]^x[362]^x[352]^x[309]^x[298]^x[74]^x[68];
	y[9]=x[383]^x[361]^x[308]^x[297]^x[73]^x[67];
	y[8]=x[382]^x[360]^x[307]^x[296]^x[72]^x[66];
	y[7]=x[381]^x[359]^x[306]^x[295]^x[71]^x[65];
	y[6]=x[380]^x[358]^x[305]^x[294]^x[70]^x[64];
	y[5]=x[379]^x[357]^x[304]^x[293]^x[138]^x[69];
	y[4]=x[378]^x[356]^x[303]^x[292]^x[137]^x[68];
	y[3]=x[377]^x[355]^x[302]^x[291]^x[136]^x[67];
	y[2]=x[376]^x[354]^x[301]^x[290]^x[135]^x[66];
	y[1]=x[375]^x[353]^x[300]^x[289]^x[134]^x[65];
	y[0]=x[374]^x[352]^x[299]^x[288]^x[133]^x[64];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint13(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[341]^x[331]^x[320]^x[287]^x[286]^x[277]^x[275]^x[266]^x[63]^x[57]^x[51]^x[45];
	y[30]=x[351]^x[350]^x[340]^x[286]^x[285]^x[276]^x[274]^x[265]^x[62]^x[56]^x[50]^x[44];
	y[29]=x[350]^x[349]^x[339]^x[285]^x[284]^x[275]^x[273]^x[264]^x[61]^x[55]^x[49]^x[43];
	y[28]=x[349]^x[348]^x[338]^x[284]^x[283]^x[274]^x[272]^x[263]^x[60]^x[54]^x[48]^x[42];
	y[27]=x[348]^x[347]^x[337]^x[283]^x[282]^x[273]^x[271]^x[262]^x[59]^x[53]^x[47]^x[41];
	y[26]=x[347]^x[346]^x[336]^x[282]^x[281]^x[272]^x[270]^x[261]^x[127]^x[106]^x[58]^x[52]^x[46]^x[40];
	y[25]=x[346]^x[345]^x[335]^x[281]^x[280]^x[271]^x[269]^x[260]^x[126]^x[105]^x[57]^x[51]^x[45]^x[39];
	y[24]=x[345]^x[344]^x[334]^x[280]^x[279]^x[270]^x[268]^x[259]^x[125]^x[104]^x[56]^x[50]^x[44]^x[38];
	y[23]=x[344]^x[343]^x[333]^x[279]^x[278]^x[269]^x[267]^x[258]^x[124]^x[103]^x[55]^x[49]^x[43]^x[37];
	y[22]=x[343]^x[342]^x[332]^x[278]^x[277]^x[268]^x[266]^x[257]^x[123]^x[102]^x[54]^x[48]^x[42]^x[36];
	y[21]=x[342]^x[341]^x[331]^x[277]^x[276]^x[267]^x[265]^x[256]^x[122]^x[101]^x[53]^x[47]^x[41]^x[35];
	y[20]=x[341]^x[340]^x[330]^x[287]^x[276]^x[275]^x[264]^x[52]^x[46]^x[40]^x[34];
	y[19]=x[340]^x[339]^x[329]^x[286]^x[275]^x[274]^x[263]^x[51]^x[45]^x[39]^x[33];
	y[18]=x[339]^x[338]^x[328]^x[285]^x[274]^x[273]^x[262]^x[50]^x[44]^x[38]^x[32];
	y[17]=x[338]^x[337]^x[327]^x[284]^x[273]^x[272]^x[261]^x[49]^x[43]^x[37];
	y[16]=x[337]^x[336]^x[326]^x[283]^x[272]^x[271]^x[260]^x[48]^x[42]^x[36];
	y[15]=x[336]^x[335]^x[325]^x[282]^x[271]^x[270]^x[259]^x[47]^x[41]^x[35];
	y[14]=x[335]^x[334]^x[324]^x[281]^x[270]^x[269]^x[258]^x[46]^x[40]^x[34];
	y[13]=x[334]^x[333]^x[323]^x[280]^x[269]^x[268]^x[257]^x[45]^x[39]^x[33];
	y[12]=x[333]^x[332]^x[322]^x[279]^x[268]^x[267]^x[256]^x[44]^x[38]^x[32];
	y[11]=x[332]^x[331]^x[321]^x[278]^x[267]^x[43]^x[37];
	y[10]=x[331]^x[330]^x[320]^x[277]^x[266]^x[42]^x[36];
	y[9]=x[351]^x[329]^x[276]^x[265]^x[41]^x[35];
	y[8]=x[350]^x[328]^x[275]^x[264]^x[40]^x[34];
	y[7]=x[349]^x[327]^x[274]^x[263]^x[39]^x[33];
	y[6]=x[348]^x[326]^x[273]^x[262]^x[38]^x[32];
	y[5]=x[347]^x[325]^x[272]^x[261]^x[106]^x[37];
	y[4]=x[346]^x[324]^x[271]^x[260]^x[105]^x[36];
	y[3]=x[345]^x[323]^x[270]^x[259]^x[104]^x[35];
	y[2]=x[344]^x[322]^x[269]^x[258]^x[103]^x[34];
	y[1]=x[343]^x[321]^x[268]^x[257]^x[102]^x[33];
	y[0]=x[342]^x[320]^x[267]^x[256]^x[101]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint14(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[319]^x[309]^x[299]^x[288]^x[255]^x[254]^x[245]^x[243]^x[234]^x[31]^x[25]^x[19]^x[13];
	y[30]=x[319]^x[318]^x[308]^x[254]^x[253]^x[244]^x[242]^x[233]^x[30]^x[24]^x[18]^x[12];
	y[29]=x[318]^x[317]^x[307]^x[253]^x[252]^x[243]^x[241]^x[232]^x[29]^x[23]^x[17]^x[11];
	y[28]=x[317]^x[316]^x[306]^x[252]^x[251]^x[242]^x[240]^x[231]^x[28]^x[22]^x[16]^x[10];
	y[27]=x[316]^x[315]^x[305]^x[251]^x[250]^x[241]^x[239]^x[230]^x[27]^x[21]^x[15]^x[9];
	y[26]=x[315]^x[314]^x[304]^x[250]^x[249]^x[240]^x[238]^x[229]^x[95]^x[74]^x[26]^x[20]^x[14]^x[8];
	y[25]=x[314]^x[313]^x[303]^x[249]^x[248]^x[239]^x[237]^x[228]^x[94]^x[73]^x[25]^x[19]^x[13]^x[7];
	y[24]=x[313]^x[312]^x[302]^x[248]^x[247]^x[238]^x[236]^x[227]^x[93]^x[72]^x[24]^x[18]^x[12]^x[6];
	y[23]=x[312]^x[311]^x[301]^x[247]^x[246]^x[237]^x[235]^x[226]^x[92]^x[71]^x[23]^x[17]^x[11]^x[5];
	y[22]=x[311]^x[310]^x[300]^x[246]^x[245]^x[236]^x[234]^x[225]^x[91]^x[70]^x[22]^x[16]^x[10]^x[4];
	y[21]=x[310]^x[309]^x[299]^x[245]^x[244]^x[235]^x[233]^x[224]^x[90]^x[69]^x[21]^x[15]^x[9]^x[3];
	y[20]=x[309]^x[308]^x[298]^x[255]^x[244]^x[243]^x[232]^x[20]^x[14]^x[8]^x[2];
	y[19]=x[308]^x[307]^x[297]^x[254]^x[243]^x[242]^x[231]^x[19]^x[13]^x[7]^x[1];
	y[18]=x[307]^x[306]^x[296]^x[253]^x[242]^x[241]^x[230]^x[18]^x[12]^x[6]^x[0];
	y[17]=x[306]^x[305]^x[295]^x[252]^x[241]^x[240]^x[229]^x[17]^x[11]^x[5];
	y[16]=x[305]^x[304]^x[294]^x[251]^x[240]^x[239]^x[228]^x[16]^x[10]^x[4];
	y[15]=x[304]^x[303]^x[293]^x[250]^x[239]^x[238]^x[227]^x[15]^x[9]^x[3];
	y[14]=x[303]^x[302]^x[292]^x[249]^x[238]^x[237]^x[226]^x[14]^x[8]^x[2];
	y[13]=x[302]^x[301]^x[291]^x[248]^x[237]^x[236]^x[225]^x[13]^x[7]^x[1];
	y[12]=x[301]^x[300]^x[290]^x[247]^x[236]^x[235]^x[224]^x[12]^x[6]^x[0];
	y[11]=x[300]^x[299]^x[289]^x[246]^x[235]^x[11]^x[5];
	y[10]=x[299]^x[298]^x[288]^x[245]^x[234]^x[10]^x[4];
	y[9]=x[319]^x[297]^x[244]^x[233]^x[9]^x[3];
	y[8]=x[318]^x[296]^x[243]^x[232]^x[8]^x[2];
	y[7]=x[317]^x[295]^x[242]^x[231]^x[7]^x[1];
	y[6]=x[316]^x[294]^x[241]^x[230]^x[6]^x[0];
	y[5]=x[315]^x[293]^x[240]^x[229]^x[74]^x[5];
	y[4]=x[314]^x[292]^x[239]^x[228]^x[73]^x[4];
	y[3]=x[313]^x[291]^x[238]^x[227]^x[72]^x[3];
	y[2]=x[312]^x[290]^x[237]^x[226]^x[71]^x[2];
	y[1]=x[311]^x[289]^x[236]^x[225]^x[70]^x[1];
	y[0]=x[310]^x[288]^x[235]^x[224]^x[69]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint15(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[377]^x[376]^x[373]^x[371]^x[367]^x[365]^x[362]^x[356]^x[287]^x[277]^x[267]^x[256]^x[223]^x[222]^x[213]^x[211]^x[202]^x[159]^x[135];
	y[30]=x[382]^x[381]^x[376]^x[375]^x[372]^x[370]^x[366]^x[364]^x[361]^x[355]^x[287]^x[286]^x[276]^x[222]^x[221]^x[212]^x[210]^x[201]^x[158]^x[134];
	y[29]=x[381]^x[380]^x[375]^x[374]^x[371]^x[369]^x[365]^x[363]^x[360]^x[354]^x[286]^x[285]^x[275]^x[221]^x[220]^x[211]^x[209]^x[200]^x[157]^x[133];
	y[28]=x[380]^x[379]^x[374]^x[373]^x[370]^x[368]^x[364]^x[362]^x[359]^x[353]^x[285]^x[284]^x[274]^x[220]^x[219]^x[210]^x[208]^x[199]^x[156]^x[132];
	y[27]=x[379]^x[378]^x[373]^x[372]^x[369]^x[367]^x[363]^x[361]^x[358]^x[352]^x[284]^x[283]^x[273]^x[219]^x[218]^x[209]^x[207]^x[198]^x[155]^x[131];
	y[26]=x[383]^x[378]^x[377]^x[372]^x[371]^x[368]^x[366]^x[360]^x[357]^x[283]^x[282]^x[272]^x[218]^x[217]^x[208]^x[206]^x[197]^x[154]^x[130]^x[63]^x[42];
	y[25]=x[382]^x[377]^x[376]^x[371]^x[370]^x[367]^x[365]^x[359]^x[356]^x[282]^x[281]^x[271]^x[217]^x[216]^x[207]^x[205]^x[196]^x[153]^x[129]^x[62]^x[41];
	y[24]=x[381]^x[376]^x[375]^x[370]^x[369]^x[366]^x[364]^x[358]^x[355]^x[281]^x[280]^x[270]^x[216]^x[215]^x[206]^x[204]^x[195]^x[152]^x[128]^x[61]^x[40];
	y[23]=x[380]^x[375]^x[374]^x[369]^x[368]^x[365]^x[363]^x[357]^x[354]^x[280]^x[279]^x[269]^x[215]^x[214]^x[205]^x[203]^x[194]^x[151]^x[60]^x[39];
	y[22]=x[379]^x[374]^x[373]^x[368]^x[367]^x[364]^x[362]^x[356]^x[353]^x[279]^x[278]^x[268]^x[214]^x[213]^x[204]^x[202]^x[193]^x[150]^x[59]^x[38];
	y[21]=x[378]^x[373]^x[372]^x[367]^x[366]^x[363]^x[361]^x[355]^x[352]^x[278]^x[277]^x[267]^x[213]^x[212]^x[203]^x[201]^x[192]^x[149]^x[58]^x[37];
	y[20]=x[383]^x[377]^x[372]^x[371]^x[366]^x[365]^x[360]^x[354]^x[277]^x[276]^x[266]^x[223]^x[212]^x[211]^x[200]^x[148];
	y[19]=x[382]^x[376]^x[371]^x[370]^x[365]^x[364]^x[359]^x[353]^x[276]^x[275]^x[265]^x[222]^x[211]^x[210]^x[199]^x[147];
	y[18]=x[381]^x[375]^x[370]^x[369]^x[364]^x[363]^x[358]^x[352]^x[275]^x[274]^x[264]^x[221]^x[210]^x[209]^x[198]^x[146];
	y[17]=x[380]^x[374]^x[369]^x[368]^x[363]^x[357]^x[274]^x[273]^x[263]^x[220]^x[209]^x[208]^x[197]^x[145];
	y[16]=x[379]^x[373]^x[368]^x[367]^x[362]^x[356]^x[273]^x[272]^x[262]^x[219]^x[208]^x[207]^x[196]^x[144];
	y[15]=x[378]^x[372]^x[367]^x[366]^x[361]^x[355]^x[272]^x[271]^x[261]^x[218]^x[207]^x[206]^x[195]^x[143];
	y[14]=x[377]^x[371]^x[366]^x[365]^x[360]^x[354]^x[271]^x[270]^x[260]^x[217]^x[206]^x[205]^x[194]^x[142];
	y[13]=x[376]^x[370]^x[365]^x[364]^x[359]^x[353]^x[270]^x[269]^x[259]^x[216]^x[205]^x[204]^x[193]^x[141];
	y[12]=x[375]^x[369]^x[364]^x[363]^x[358]^x[352]^x[269]^x[268]^x[258]^x[215]^x[204]^x[203]^x[192]^x[140];
	y[11]=x[374]^x[368]^x[363]^x[357]^x[268]^x[267]^x[257]^x[214]^x[203]^x[139];
	y[10]=x[373]^x[367]^x[362]^x[356]^x[267]^x[266]^x[256]^x[213]^x[202]^x[138];
	y[9]=x[372]^x[366]^x[361]^x[355]^x[287]^x[265]^x[212]^x[201]^x[137];
	y[8]=x[371]^x[365]^x[360]^x[354]^x[286]^x[264]^x[211]^x[200]^x[136];
	y[7]=x[370]^x[364]^x[359]^x[353]^x[285]^x[263]^x[210]^x[199]^x[135];
	y[6]=x[369]^x[363]^x[358]^x[352]^x[284]^x[262]^x[209]^x[198]^x[134];
	y[5]=x[368]^x[357]^x[283]^x[261]^x[208]^x[197]^x[133]^x[42];
	y[4]=x[367]^x[356]^x[282]^x[260]^x[207]^x[196]^x[132]^x[41];
	y[3]=x[366]^x[355]^x[281]^x[259]^x[206]^x[195]^x[131]^x[40];
	y[2]=x[365]^x[354]^x[280]^x[258]^x[205]^x[194]^x[130]^x[39];
	y[1]=x[364]^x[353]^x[279]^x[257]^x[204]^x[193]^x[129]^x[38];
	y[0]=x[363]^x[352]^x[278]^x[256]^x[203]^x[192]^x[128]^x[37];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint16(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[350]^x[345]^x[344]^x[341]^x[339]^x[335]^x[333]^x[330]^x[324]^x[255]^x[245]^x[235]^x[224]^x[191]^x[190]^x[181]^x[179]^x[170]^x[127]^x[103];
	y[30]=x[350]^x[349]^x[344]^x[343]^x[340]^x[338]^x[334]^x[332]^x[329]^x[323]^x[255]^x[254]^x[244]^x[190]^x[189]^x[180]^x[178]^x[169]^x[126]^x[102];
	y[29]=x[349]^x[348]^x[343]^x[342]^x[339]^x[337]^x[333]^x[331]^x[328]^x[322]^x[254]^x[253]^x[243]^x[189]^x[188]^x[179]^x[177]^x[168]^x[125]^x[101];
	y[28]=x[348]^x[347]^x[342]^x[341]^x[338]^x[336]^x[332]^x[330]^x[327]^x[321]^x[253]^x[252]^x[242]^x[188]^x[187]^x[178]^x[176]^x[167]^x[124]^x[100];
	y[27]=x[347]^x[346]^x[341]^x[340]^x[337]^x[335]^x[331]^x[329]^x[326]^x[320]^x[252]^x[251]^x[241]^x[187]^x[186]^x[177]^x[175]^x[166]^x[123]^x[99];
	y[26]=x[351]^x[346]^x[345]^x[340]^x[339]^x[336]^x[334]^x[328]^x[325]^x[251]^x[250]^x[240]^x[186]^x[185]^x[176]^x[174]^x[165]^x[122]^x[98]^x[31]^x[10];
	y[25]=x[350]^x[345]^x[344]^x[339]^x[338]^x[335]^x[333]^x[327]^x[324]^x[250]^x[249]^x[239]^x[185]^x[184]^x[175]^x[173]^x[164]^x[121]^x[97]^x[30]^x[9];
	y[24]=x[349]^x[344]^x[343]^x[338]^x[337]^x[334]^x[332]^x[326]^x[323]^x[249]^x[248]^x[238]^x[184]^x[183]^x[174]^x[172]^x[163]^x[120]^x[96]^x[29]^x[8];
	y[23]=x[348]^x[343]^x[342]^x[337]^x[336]^x[333]^x[331]^x[325]^x[322]^x[248]^x[247]^x[237]^x[183]^x[182]^x[173]^x[171]^x[162]^x[119]^x[28]^x[7];
	y[22]=x[347]^x[342]^x[341]^x[336]^x[335]^x[332]^x[330]^x[324]^x[321]^x[247]^x[246]^x[236]^x[182]^x[181]^x[172]^x[170]^x[161]^x[118]^x[27]^x[6];
	y[21]=x[346]^x[341]^x[340]^x[335]^x[334]^x[331]^x[329]^x[323]^x[320]^x[246]^x[245]^x[235]^x[181]^x[180]^x[171]^x[169]^x[160]^x[117]^x[26]^x[5];
	y[20]=x[351]^x[345]^x[340]^x[339]^x[334]^x[333]^x[328]^x[322]^x[245]^x[244]^x[234]^x[191]^x[180]^x[179]^x[168]^x[116];
	y[19]=x[350]^x[344]^x[339]^x[338]^x[333]^x[332]^x[327]^x[321]^x[244]^x[243]^x[233]^x[190]^x[179]^x[178]^x[167]^x[115];
	y[18]=x[349]^x[343]^x[338]^x[337]^x[332]^x[331]^x[326]^x[320]^x[243]^x[242]^x[232]^x[189]^x[178]^x[177]^x[166]^x[114];
	y[17]=x[348]^x[342]^x[337]^x[336]^x[331]^x[325]^x[242]^x[241]^x[231]^x[188]^x[177]^x[176]^x[165]^x[113];
	y[16]=x[347]^x[341]^x[336]^x[335]^x[330]^x[324]^x[241]^x[240]^x[230]^x[187]^x[176]^x[175]^x[164]^x[112];
	y[15]=x[346]^x[340]^x[335]^x[334]^x[329]^x[323]^x[240]^x[239]^x[229]^x[186]^x[175]^x[174]^x[163]^x[111];
	y[14]=x[345]^x[339]^x[334]^x[333]^x[328]^x[322]^x[239]^x[238]^x[228]^x[185]^x[174]^x[173]^x[162]^x[110];
	y[13]=x[344]^x[338]^x[333]^x[332]^x[327]^x[321]^x[238]^x[237]^x[227]^x[184]^x[173]^x[172]^x[161]^x[109];
	y[12]=x[343]^x[337]^x[332]^x[331]^x[326]^x[320]^x[237]^x[236]^x[226]^x[183]^x[172]^x[171]^x[160]^x[108];
	y[11]=x[342]^x[336]^x[331]^x[325]^x[236]^x[235]^x[225]^x[182]^x[171]^x[107];
	y[10]=x[341]^x[335]^x[330]^x[324]^x[235]^x[234]^x[224]^x[181]^x[170]^x[106];
	y[9]=x[340]^x[334]^x[329]^x[323]^x[255]^x[233]^x[180]^x[169]^x[105];
	y[8]=x[339]^x[333]^x[328]^x[322]^x[254]^x[232]^x[179]^x[168]^x[104];
	y[7]=x[338]^x[332]^x[327]^x[321]^x[253]^x[231]^x[178]^x[167]^x[103];
	y[6]=x[337]^x[331]^x[326]^x[320]^x[252]^x[230]^x[177]^x[166]^x[102];
	y[5]=x[336]^x[325]^x[251]^x[229]^x[176]^x[165]^x[101]^x[10];
	y[4]=x[335]^x[324]^x[250]^x[228]^x[175]^x[164]^x[100]^x[9];
	y[3]=x[334]^x[323]^x[249]^x[227]^x[174]^x[163]^x[99]^x[8];
	y[2]=x[333]^x[322]^x[248]^x[226]^x[173]^x[162]^x[98]^x[7];
	y[1]=x[332]^x[321]^x[247]^x[225]^x[172]^x[161]^x[97]^x[6];
	y[0]=x[331]^x[320]^x[246]^x[224]^x[171]^x[160]^x[96]^x[5];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint17(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[319]^x[318]^x[313]^x[312]^x[309]^x[307]^x[303]^x[301]^x[298]^x[292]^x[223]^x[213]^x[203]^x[192]^x[159]^x[158]^x[149]^x[147]^x[138]^x[95]^x[71];
	y[30]=x[318]^x[317]^x[312]^x[311]^x[308]^x[306]^x[302]^x[300]^x[297]^x[291]^x[223]^x[222]^x[212]^x[158]^x[157]^x[148]^x[146]^x[137]^x[94]^x[70];
	y[29]=x[317]^x[316]^x[311]^x[310]^x[307]^x[305]^x[301]^x[299]^x[296]^x[290]^x[222]^x[221]^x[211]^x[157]^x[156]^x[147]^x[145]^x[136]^x[93]^x[69];
	y[28]=x[316]^x[315]^x[310]^x[309]^x[306]^x[304]^x[300]^x[298]^x[295]^x[289]^x[221]^x[220]^x[210]^x[156]^x[155]^x[146]^x[144]^x[135]^x[92]^x[68];
	y[27]=x[315]^x[314]^x[309]^x[308]^x[305]^x[303]^x[299]^x[297]^x[294]^x[288]^x[220]^x[219]^x[209]^x[155]^x[154]^x[145]^x[143]^x[134]^x[91]^x[67];
	y[26]=x[383]^x[319]^x[314]^x[313]^x[308]^x[307]^x[304]^x[302]^x[296]^x[293]^x[219]^x[218]^x[208]^x[159]^x[154]^x[144]^x[142]^x[138]^x[133]^x[132]^x[90]^x[66];
	y[25]=x[382]^x[318]^x[313]^x[312]^x[307]^x[306]^x[303]^x[301]^x[295]^x[292]^x[218]^x[217]^x[207]^x[158]^x[153]^x[143]^x[141]^x[137]^x[132]^x[131]^x[89]^x[65];
	y[24]=x[381]^x[317]^x[312]^x[311]^x[306]^x[305]^x[302]^x[300]^x[294]^x[291]^x[217]^x[216]^x[206]^x[157]^x[152]^x[142]^x[140]^x[136]^x[131]^x[130]^x[88]^x[64];
	y[23]=x[380]^x[316]^x[311]^x[310]^x[305]^x[304]^x[301]^x[299]^x[293]^x[290]^x[216]^x[215]^x[205]^x[156]^x[151]^x[141]^x[139]^x[135]^x[130]^x[129]^x[87];
	y[22]=x[379]^x[315]^x[310]^x[309]^x[304]^x[303]^x[300]^x[298]^x[292]^x[289]^x[215]^x[214]^x[204]^x[155]^x[150]^x[140]^x[138]^x[134]^x[129]^x[128]^x[86];
	y[21]=x[378]^x[314]^x[309]^x[308]^x[303]^x[302]^x[299]^x[297]^x[291]^x[288]^x[214]^x[213]^x[203]^x[154]^x[149]^x[139]^x[137]^x[133]^x[128]^x[85];
	y[20]=x[319]^x[313]^x[308]^x[307]^x[302]^x[301]^x[296]^x[290]^x[213]^x[212]^x[202]^x[159]^x[148]^x[147]^x[136]^x[84];
	y[19]=x[318]^x[312]^x[307]^x[306]^x[301]^x[300]^x[295]^x[289]^x[212]^x[211]^x[201]^x[158]^x[147]^x[146]^x[135]^x[83];
	y[18]=x[317]^x[311]^x[306]^x[305]^x[300]^x[299]^x[294]^x[288]^x[211]^x[210]^x[200]^x[157]^x[146]^x[145]^x[134]^x[82];
	y[17]=x[316]^x[310]^x[305]^x[304]^x[299]^x[293]^x[210]^x[209]^x[199]^x[156]^x[145]^x[144]^x[133]^x[81];
	y[16]=x[315]^x[309]^x[304]^x[303]^x[298]^x[292]^x[209]^x[208]^x[198]^x[155]^x[144]^x[143]^x[132]^x[80];
	y[15]=x[314]^x[308]^x[303]^x[302]^x[297]^x[291]^x[208]^x[207]^x[197]^x[154]^x[143]^x[142]^x[131]^x[79];
	y[14]=x[313]^x[307]^x[302]^x[301]^x[296]^x[290]^x[207]^x[206]^x[196]^x[153]^x[142]^x[141]^x[130]^x[78];
	y[13]=x[312]^x[306]^x[301]^x[300]^x[295]^x[289]^x[206]^x[205]^x[195]^x[152]^x[141]^x[140]^x[129]^x[77];
	y[12]=x[311]^x[305]^x[300]^x[299]^x[294]^x[288]^x[205]^x[204]^x[194]^x[151]^x[140]^x[139]^x[128]^x[76];
	y[11]=x[310]^x[304]^x[299]^x[293]^x[204]^x[203]^x[193]^x[150]^x[139]^x[75];
	y[10]=x[309]^x[303]^x[298]^x[292]^x[203]^x[202]^x[192]^x[149]^x[138]^x[74];
	y[9]=x[308]^x[302]^x[297]^x[291]^x[223]^x[201]^x[148]^x[137]^x[73];
	y[8]=x[307]^x[301]^x[296]^x[290]^x[222]^x[200]^x[147]^x[136]^x[72];
	y[7]=x[306]^x[300]^x[295]^x[289]^x[221]^x[199]^x[146]^x[135]^x[71];
	y[6]=x[305]^x[299]^x[294]^x[288]^x[220]^x[198]^x[145]^x[134]^x[70];
	y[5]=x[373]^x[362]^x[304]^x[293]^x[219]^x[197]^x[144]^x[138]^x[133]^x[132]^x[69];
	y[4]=x[372]^x[361]^x[303]^x[292]^x[218]^x[196]^x[143]^x[137]^x[132]^x[131]^x[68];
	y[3]=x[371]^x[360]^x[302]^x[291]^x[217]^x[195]^x[142]^x[136]^x[131]^x[130]^x[67];
	y[2]=x[370]^x[359]^x[301]^x[290]^x[216]^x[194]^x[141]^x[135]^x[130]^x[129]^x[66];
	y[1]=x[369]^x[358]^x[300]^x[289]^x[215]^x[193]^x[140]^x[134]^x[129]^x[128]^x[65];
	y[0]=x[368]^x[357]^x[299]^x[288]^x[214]^x[192]^x[139]^x[133]^x[128]^x[64];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint18(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[287]^x[286]^x[281]^x[280]^x[277]^x[275]^x[271]^x[269]^x[266]^x[260]^x[191]^x[181]^x[171]^x[160]^x[127]^x[126]^x[117]^x[115]^x[106]^x[63]^x[39];
	y[30]=x[286]^x[285]^x[280]^x[279]^x[276]^x[274]^x[270]^x[268]^x[265]^x[259]^x[191]^x[190]^x[180]^x[126]^x[125]^x[116]^x[114]^x[105]^x[62]^x[38];
	y[29]=x[285]^x[284]^x[279]^x[278]^x[275]^x[273]^x[269]^x[267]^x[264]^x[258]^x[190]^x[189]^x[179]^x[125]^x[124]^x[115]^x[113]^x[104]^x[61]^x[37];
	y[28]=x[284]^x[283]^x[278]^x[277]^x[274]^x[272]^x[268]^x[266]^x[263]^x[257]^x[189]^x[188]^x[178]^x[124]^x[123]^x[114]^x[112]^x[103]^x[60]^x[36];
	y[27]=x[283]^x[282]^x[277]^x[276]^x[273]^x[271]^x[267]^x[265]^x[262]^x[256]^x[188]^x[187]^x[177]^x[123]^x[122]^x[113]^x[111]^x[102]^x[59]^x[35];
	y[26]=x[351]^x[287]^x[282]^x[281]^x[276]^x[275]^x[272]^x[270]^x[264]^x[261]^x[187]^x[186]^x[176]^x[127]^x[122]^x[112]^x[110]^x[106]^x[101]^x[100]^x[58]^x[34];
	y[25]=x[350]^x[286]^x[281]^x[280]^x[275]^x[274]^x[271]^x[269]^x[263]^x[260]^x[186]^x[185]^x[175]^x[126]^x[121]^x[111]^x[109]^x[105]^x[100]^x[99]^x[57]^x[33];
	y[24]=x[349]^x[285]^x[280]^x[279]^x[274]^x[273]^x[270]^x[268]^x[262]^x[259]^x[185]^x[184]^x[174]^x[125]^x[120]^x[110]^x[108]^x[104]^x[99]^x[98]^x[56]^x[32];
	y[23]=x[348]^x[284]^x[279]^x[278]^x[273]^x[272]^x[269]^x[267]^x[261]^x[258]^x[184]^x[183]^x[173]^x[124]^x[119]^x[109]^x[107]^x[103]^x[98]^x[97]^x[55];
	y[22]=x[347]^x[283]^x[278]^x[277]^x[272]^x[271]^x[268]^x[266]^x[260]^x[257]^x[183]^x[182]^x[172]^x[123]^x[118]^x[108]^x[106]^x[102]^x[97]^x[96]^x[54];
	y[21]=x[346]^x[282]^x[277]^x[276]^x[271]^x[270]^x[267]^x[265]^x[259]^x[256]^x[182]^x[181]^x[171]^x[122]^x[117]^x[107]^x[105]^x[101]^x[96]^x[53];
	y[20]=x[287]^x[281]^x[276]^x[275]^x[270]^x[269]^x[264]^x[258]^x[181]^x[180]^x[170]^x[127]^x[116]^x[115]^x[104]^x[52];
	y[19]=x[286]^x[280]^x[275]^x[274]^x[269]^x[268]^x[263]^x[257]^x[180]^x[179]^x[169]^x[126]^x[115]^x[114]^x[103]^x[51];
	y[18]=x[285]^x[279]^x[274]^x[273]^x[268]^x[267]^x[262]^x[256]^x[179]^x[178]^x[168]^x[125]^x[114]^x[113]^x[102]^x[50];
	y[17]=x[284]^x[278]^x[273]^x[272]^x[267]^x[261]^x[178]^x[177]^x[167]^x[124]^x[113]^x[112]^x[101]^x[49];
	y[16]=x[283]^x[277]^x[272]^x[271]^x[266]^x[260]^x[177]^x[176]^x[166]^x[123]^x[112]^x[111]^x[100]^x[48];
	y[15]=x[282]^x[276]^x[271]^x[270]^x[265]^x[259]^x[176]^x[175]^x[165]^x[122]^x[111]^x[110]^x[99]^x[47];
	y[14]=x[281]^x[275]^x[270]^x[269]^x[264]^x[258]^x[175]^x[174]^x[164]^x[121]^x[110]^x[109]^x[98]^x[46];
	y[13]=x[280]^x[274]^x[269]^x[268]^x[263]^x[257]^x[174]^x[173]^x[163]^x[120]^x[109]^x[108]^x[97]^x[45];
	y[12]=x[279]^x[273]^x[268]^x[267]^x[262]^x[256]^x[173]^x[172]^x[162]^x[119]^x[108]^x[107]^x[96]^x[44];
	y[11]=x[278]^x[272]^x[267]^x[261]^x[172]^x[171]^x[161]^x[118]^x[107]^x[43];
	y[10]=x[277]^x[271]^x[266]^x[260]^x[171]^x[170]^x[160]^x[117]^x[106]^x[42];
	y[9]=x[276]^x[270]^x[265]^x[259]^x[191]^x[169]^x[116]^x[105]^x[41];
	y[8]=x[275]^x[269]^x[264]^x[258]^x[190]^x[168]^x[115]^x[104]^x[40];
	y[7]=x[274]^x[268]^x[263]^x[257]^x[189]^x[167]^x[114]^x[103]^x[39];
	y[6]=x[273]^x[267]^x[262]^x[256]^x[188]^x[166]^x[113]^x[102]^x[38];
	y[5]=x[341]^x[330]^x[272]^x[261]^x[187]^x[165]^x[112]^x[106]^x[101]^x[100]^x[37];
	y[4]=x[340]^x[329]^x[271]^x[260]^x[186]^x[164]^x[111]^x[105]^x[100]^x[99]^x[36];
	y[3]=x[339]^x[328]^x[270]^x[259]^x[185]^x[163]^x[110]^x[104]^x[99]^x[98]^x[35];
	y[2]=x[338]^x[327]^x[269]^x[258]^x[184]^x[162]^x[109]^x[103]^x[98]^x[97]^x[34];
	y[1]=x[337]^x[326]^x[268]^x[257]^x[183]^x[161]^x[108]^x[102]^x[97]^x[96]^x[33];
	y[0]=x[336]^x[325]^x[267]^x[256]^x[182]^x[160]^x[107]^x[101]^x[96]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint19(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[255]^x[254]^x[249]^x[248]^x[245]^x[243]^x[239]^x[237]^x[234]^x[228]^x[159]^x[149]^x[139]^x[128]^x[95]^x[94]^x[85]^x[83]^x[74]^x[31]^x[7];
	y[30]=x[254]^x[253]^x[248]^x[247]^x[244]^x[242]^x[238]^x[236]^x[233]^x[227]^x[159]^x[158]^x[148]^x[94]^x[93]^x[84]^x[82]^x[73]^x[30]^x[6];
	y[29]=x[253]^x[252]^x[247]^x[246]^x[243]^x[241]^x[237]^x[235]^x[232]^x[226]^x[158]^x[157]^x[147]^x[93]^x[92]^x[83]^x[81]^x[72]^x[29]^x[5];
	y[28]=x[252]^x[251]^x[246]^x[245]^x[242]^x[240]^x[236]^x[234]^x[231]^x[225]^x[157]^x[156]^x[146]^x[92]^x[91]^x[82]^x[80]^x[71]^x[28]^x[4];
	y[27]=x[251]^x[250]^x[245]^x[244]^x[241]^x[239]^x[235]^x[233]^x[230]^x[224]^x[156]^x[155]^x[145]^x[91]^x[90]^x[81]^x[79]^x[70]^x[27]^x[3];
	y[26]=x[319]^x[255]^x[250]^x[249]^x[244]^x[243]^x[240]^x[238]^x[232]^x[229]^x[155]^x[154]^x[144]^x[95]^x[90]^x[80]^x[78]^x[74]^x[69]^x[68]^x[26]^x[2];
	y[25]=x[318]^x[254]^x[249]^x[248]^x[243]^x[242]^x[239]^x[237]^x[231]^x[228]^x[154]^x[153]^x[143]^x[94]^x[89]^x[79]^x[77]^x[73]^x[68]^x[67]^x[25]^x[1];
	y[24]=x[317]^x[253]^x[248]^x[247]^x[242]^x[241]^x[238]^x[236]^x[230]^x[227]^x[153]^x[152]^x[142]^x[93]^x[88]^x[78]^x[76]^x[72]^x[67]^x[66]^x[24]^x[0];
	y[23]=x[316]^x[252]^x[247]^x[246]^x[241]^x[240]^x[237]^x[235]^x[229]^x[226]^x[152]^x[151]^x[141]^x[92]^x[87]^x[77]^x[75]^x[71]^x[66]^x[65]^x[23];
	y[22]=x[315]^x[251]^x[246]^x[245]^x[240]^x[239]^x[236]^x[234]^x[228]^x[225]^x[151]^x[150]^x[140]^x[91]^x[86]^x[76]^x[74]^x[70]^x[65]^x[64]^x[22];
	y[21]=x[314]^x[250]^x[245]^x[244]^x[239]^x[238]^x[235]^x[233]^x[227]^x[224]^x[150]^x[149]^x[139]^x[90]^x[85]^x[75]^x[73]^x[69]^x[64]^x[21];
	y[20]=x[255]^x[249]^x[244]^x[243]^x[238]^x[237]^x[232]^x[226]^x[149]^x[148]^x[138]^x[95]^x[84]^x[83]^x[72]^x[20];
	y[19]=x[254]^x[248]^x[243]^x[242]^x[237]^x[236]^x[231]^x[225]^x[148]^x[147]^x[137]^x[94]^x[83]^x[82]^x[71]^x[19];
	y[18]=x[253]^x[247]^x[242]^x[241]^x[236]^x[235]^x[230]^x[224]^x[147]^x[146]^x[136]^x[93]^x[82]^x[81]^x[70]^x[18];
	y[17]=x[252]^x[246]^x[241]^x[240]^x[235]^x[229]^x[146]^x[145]^x[135]^x[92]^x[81]^x[80]^x[69]^x[17];
	y[16]=x[251]^x[245]^x[240]^x[239]^x[234]^x[228]^x[145]^x[144]^x[134]^x[91]^x[80]^x[79]^x[68]^x[16];
	y[15]=x[250]^x[244]^x[239]^x[238]^x[233]^x[227]^x[144]^x[143]^x[133]^x[90]^x[79]^x[78]^x[67]^x[15];
	y[14]=x[249]^x[243]^x[238]^x[237]^x[232]^x[226]^x[143]^x[142]^x[132]^x[89]^x[78]^x[77]^x[66]^x[14];
	y[13]=x[248]^x[242]^x[237]^x[236]^x[231]^x[225]^x[142]^x[141]^x[131]^x[88]^x[77]^x[76]^x[65]^x[13];
	y[12]=x[247]^x[241]^x[236]^x[235]^x[230]^x[224]^x[141]^x[140]^x[130]^x[87]^x[76]^x[75]^x[64]^x[12];
	y[11]=x[246]^x[240]^x[235]^x[229]^x[140]^x[139]^x[129]^x[86]^x[75]^x[11];
	y[10]=x[245]^x[239]^x[234]^x[228]^x[139]^x[138]^x[128]^x[85]^x[74]^x[10];
	y[9]=x[244]^x[238]^x[233]^x[227]^x[159]^x[137]^x[84]^x[73]^x[9];
	y[8]=x[243]^x[237]^x[232]^x[226]^x[158]^x[136]^x[83]^x[72]^x[8];
	y[7]=x[242]^x[236]^x[231]^x[225]^x[157]^x[135]^x[82]^x[71]^x[7];
	y[6]=x[241]^x[235]^x[230]^x[224]^x[156]^x[134]^x[81]^x[70]^x[6];
	y[5]=x[309]^x[298]^x[240]^x[229]^x[155]^x[133]^x[80]^x[74]^x[69]^x[68]^x[5];
	y[4]=x[308]^x[297]^x[239]^x[228]^x[154]^x[132]^x[79]^x[73]^x[68]^x[67]^x[4];
	y[3]=x[307]^x[296]^x[238]^x[227]^x[153]^x[131]^x[78]^x[72]^x[67]^x[66]^x[3];
	y[2]=x[306]^x[295]^x[237]^x[226]^x[152]^x[130]^x[77]^x[71]^x[66]^x[65]^x[2];
	y[1]=x[305]^x[294]^x[236]^x[225]^x[151]^x[129]^x[76]^x[70]^x[65]^x[64]^x[1];
	y[0]=x[304]^x[293]^x[235]^x[224]^x[150]^x[128]^x[75]^x[69]^x[64]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint20(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[373]^x[370]^x[362]^x[359]^x[223]^x[222]^x[217]^x[216]^x[213]^x[211]^x[207]^x[205]^x[202]^x[196]^x[159]^x[153]^x[135]^x[129]^x[127]^x[117]^x[107]^x[96]^x[63]^x[62]^x[53]^x[51]^x[42];
	y[30]=x[382]^x[372]^x[369]^x[361]^x[358]^x[222]^x[221]^x[216]^x[215]^x[212]^x[210]^x[206]^x[204]^x[201]^x[195]^x[158]^x[152]^x[134]^x[128]^x[127]^x[126]^x[116]^x[62]^x[61]^x[52]^x[50]^x[41];
	y[29]=x[381]^x[371]^x[368]^x[360]^x[357]^x[221]^x[220]^x[215]^x[214]^x[211]^x[209]^x[205]^x[203]^x[200]^x[194]^x[157]^x[151]^x[133]^x[126]^x[125]^x[115]^x[61]^x[60]^x[51]^x[49]^x[40];
	y[28]=x[380]^x[370]^x[367]^x[359]^x[356]^x[220]^x[219]^x[214]^x[213]^x[210]^x[208]^x[204]^x[202]^x[199]^x[193]^x[156]^x[150]^x[132]^x[125]^x[124]^x[114]^x[60]^x[59]^x[50]^x[48]^x[39];
	y[27]=x[379]^x[369]^x[366]^x[358]^x[355]^x[219]^x[218]^x[213]^x[212]^x[209]^x[207]^x[203]^x[201]^x[198]^x[192]^x[155]^x[149]^x[131]^x[124]^x[123]^x[113]^x[59]^x[58]^x[49]^x[47]^x[38];
	y[26]=x[378]^x[368]^x[365]^x[357]^x[354]^x[287]^x[223]^x[218]^x[217]^x[212]^x[211]^x[208]^x[206]^x[200]^x[197]^x[154]^x[148]^x[130]^x[123]^x[122]^x[112]^x[63]^x[58]^x[48]^x[46]^x[42]^x[37]^x[36];
	y[25]=x[377]^x[367]^x[364]^x[356]^x[353]^x[286]^x[222]^x[217]^x[216]^x[211]^x[210]^x[207]^x[205]^x[199]^x[196]^x[153]^x[147]^x[129]^x[122]^x[121]^x[111]^x[62]^x[57]^x[47]^x[45]^x[41]^x[36]^x[35];
	y[24]=x[376]^x[366]^x[363]^x[355]^x[352]^x[285]^x[221]^x[216]^x[215]^x[210]^x[209]^x[206]^x[204]^x[198]^x[195]^x[152]^x[146]^x[128]^x[121]^x[120]^x[110]^x[61]^x[56]^x[46]^x[44]^x[40]^x[35]^x[34];
	y[23]=x[375]^x[365]^x[354]^x[284]^x[220]^x[215]^x[214]^x[209]^x[208]^x[205]^x[203]^x[197]^x[194]^x[151]^x[145]^x[120]^x[119]^x[109]^x[60]^x[55]^x[45]^x[43]^x[39]^x[34]^x[33];
	y[22]=x[374]^x[364]^x[353]^x[283]^x[219]^x[214]^x[213]^x[208]^x[207]^x[204]^x[202]^x[196]^x[193]^x[150]^x[144]^x[119]^x[118]^x[108]^x[59]^x[54]^x[44]^x[42]^x[38]^x[33]^x[32];
	y[21]=x[373]^x[363]^x[352]^x[282]^x[218]^x[213]^x[212]^x[207]^x[206]^x[203]^x[201]^x[195]^x[192]^x[149]^x[143]^x[118]^x[117]^x[107]^x[58]^x[53]^x[43]^x[41]^x[37]^x[32];
	y[20]=x[383]^x[372]^x[223]^x[217]^x[212]^x[211]^x[206]^x[205]^x[200]^x[194]^x[148]^x[142]^x[117]^x[116]^x[106]^x[63]^x[52]^x[51]^x[40];
	y[19]=x[382]^x[371]^x[222]^x[216]^x[211]^x[210]^x[205]^x[204]^x[199]^x[193]^x[147]^x[141]^x[116]^x[115]^x[105]^x[62]^x[51]^x[50]^x[39];
	y[18]=x[381]^x[370]^x[221]^x[215]^x[210]^x[209]^x[204]^x[203]^x[198]^x[192]^x[146]^x[140]^x[115]^x[114]^x[104]^x[61]^x[50]^x[49]^x[38];
	y[17]=x[380]^x[369]^x[220]^x[214]^x[209]^x[208]^x[203]^x[197]^x[145]^x[139]^x[114]^x[113]^x[103]^x[60]^x[49]^x[48]^x[37];
	y[16]=x[379]^x[368]^x[219]^x[213]^x[208]^x[207]^x[202]^x[196]^x[144]^x[138]^x[113]^x[112]^x[102]^x[59]^x[48]^x[47]^x[36];
	y[15]=x[378]^x[367]^x[218]^x[212]^x[207]^x[206]^x[201]^x[195]^x[143]^x[137]^x[112]^x[111]^x[101]^x[58]^x[47]^x[46]^x[35];
	y[14]=x[377]^x[366]^x[217]^x[211]^x[206]^x[205]^x[200]^x[194]^x[142]^x[136]^x[111]^x[110]^x[100]^x[57]^x[46]^x[45]^x[34];
	y[13]=x[376]^x[365]^x[216]^x[210]^x[205]^x[204]^x[199]^x[193]^x[141]^x[135]^x[110]^x[109]^x[99]^x[56]^x[45]^x[44]^x[33];
	y[12]=x[375]^x[364]^x[215]^x[209]^x[204]^x[203]^x[198]^x[192]^x[140]^x[134]^x[109]^x[108]^x[98]^x[55]^x[44]^x[43]^x[32];
	y[11]=x[374]^x[363]^x[214]^x[208]^x[203]^x[197]^x[139]^x[133]^x[108]^x[107]^x[97]^x[54]^x[43];
	y[10]=x[373]^x[362]^x[213]^x[207]^x[202]^x[196]^x[138]^x[132]^x[107]^x[106]^x[96]^x[53]^x[42];
	y[9]=x[372]^x[361]^x[212]^x[206]^x[201]^x[195]^x[137]^x[131]^x[127]^x[105]^x[52]^x[41];
	y[8]=x[371]^x[360]^x[211]^x[205]^x[200]^x[194]^x[136]^x[130]^x[126]^x[104]^x[51]^x[40];
	y[7]=x[370]^x[359]^x[210]^x[204]^x[199]^x[193]^x[135]^x[129]^x[125]^x[103]^x[50]^x[39];
	y[6]=x[369]^x[358]^x[209]^x[203]^x[198]^x[192]^x[134]^x[128]^x[124]^x[102]^x[49]^x[38];
	y[5]=x[368]^x[357]^x[277]^x[266]^x[208]^x[197]^x[133]^x[123]^x[101]^x[48]^x[42]^x[37]^x[36];
	y[4]=x[367]^x[356]^x[276]^x[265]^x[207]^x[196]^x[132]^x[122]^x[100]^x[47]^x[41]^x[36]^x[35];
	y[3]=x[366]^x[355]^x[275]^x[264]^x[206]^x[195]^x[131]^x[121]^x[99]^x[46]^x[40]^x[35]^x[34];
	y[2]=x[365]^x[354]^x[274]^x[263]^x[205]^x[194]^x[130]^x[120]^x[98]^x[45]^x[39]^x[34]^x[33];
	y[1]=x[364]^x[353]^x[273]^x[262]^x[204]^x[193]^x[129]^x[119]^x[97]^x[44]^x[38]^x[33]^x[32];
	y[0]=x[363]^x[352]^x[272]^x[261]^x[203]^x[192]^x[128]^x[118]^x[96]^x[43]^x[37]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint21(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[341]^x[338]^x[330]^x[327]^x[191]^x[190]^x[185]^x[184]^x[181]^x[179]^x[175]^x[173]^x[170]^x[164]^x[127]^x[121]^x[103]^x[97]^x[95]^x[85]^x[75]^x[64]^x[31]^x[30]^x[21]^x[19]^x[10];
	y[30]=x[350]^x[340]^x[337]^x[329]^x[326]^x[190]^x[189]^x[184]^x[183]^x[180]^x[178]^x[174]^x[172]^x[169]^x[163]^x[126]^x[120]^x[102]^x[96]^x[95]^x[94]^x[84]^x[30]^x[29]^x[20]^x[18]^x[9];
	y[29]=x[349]^x[339]^x[336]^x[328]^x[325]^x[189]^x[188]^x[183]^x[182]^x[179]^x[177]^x[173]^x[171]^x[168]^x[162]^x[125]^x[119]^x[101]^x[94]^x[93]^x[83]^x[29]^x[28]^x[19]^x[17]^x[8];
	y[28]=x[348]^x[338]^x[335]^x[327]^x[324]^x[188]^x[187]^x[182]^x[181]^x[178]^x[176]^x[172]^x[170]^x[167]^x[161]^x[124]^x[118]^x[100]^x[93]^x[92]^x[82]^x[28]^x[27]^x[18]^x[16]^x[7];
	y[27]=x[347]^x[337]^x[334]^x[326]^x[323]^x[187]^x[186]^x[181]^x[180]^x[177]^x[175]^x[171]^x[169]^x[166]^x[160]^x[123]^x[117]^x[99]^x[92]^x[91]^x[81]^x[27]^x[26]^x[17]^x[15]^x[6];
	y[26]=x[346]^x[336]^x[333]^x[325]^x[322]^x[255]^x[191]^x[186]^x[185]^x[180]^x[179]^x[176]^x[174]^x[168]^x[165]^x[122]^x[116]^x[98]^x[91]^x[90]^x[80]^x[31]^x[26]^x[16]^x[14]^x[10]^x[5]^x[4];
	y[25]=x[345]^x[335]^x[332]^x[324]^x[321]^x[254]^x[190]^x[185]^x[184]^x[179]^x[178]^x[175]^x[173]^x[167]^x[164]^x[121]^x[115]^x[97]^x[90]^x[89]^x[79]^x[30]^x[25]^x[15]^x[13]^x[9]^x[4]^x[3];
	y[24]=x[344]^x[334]^x[331]^x[323]^x[320]^x[253]^x[189]^x[184]^x[183]^x[178]^x[177]^x[174]^x[172]^x[166]^x[163]^x[120]^x[114]^x[96]^x[89]^x[88]^x[78]^x[29]^x[24]^x[14]^x[12]^x[8]^x[3]^x[2];
	y[23]=x[343]^x[333]^x[322]^x[252]^x[188]^x[183]^x[182]^x[177]^x[176]^x[173]^x[171]^x[165]^x[162]^x[119]^x[113]^x[88]^x[87]^x[77]^x[28]^x[23]^x[13]^x[11]^x[7]^x[2]^x[1];
	y[22]=x[342]^x[332]^x[321]^x[251]^x[187]^x[182]^x[181]^x[176]^x[175]^x[172]^x[170]^x[164]^x[161]^x[118]^x[112]^x[87]^x[86]^x[76]^x[27]^x[22]^x[12]^x[10]^x[6]^x[1]^x[0];
	y[21]=x[341]^x[331]^x[320]^x[250]^x[186]^x[181]^x[180]^x[175]^x[174]^x[171]^x[169]^x[163]^x[160]^x[117]^x[111]^x[86]^x[85]^x[75]^x[26]^x[21]^x[11]^x[9]^x[5]^x[0];
	y[20]=x[351]^x[340]^x[191]^x[185]^x[180]^x[179]^x[174]^x[173]^x[168]^x[162]^x[116]^x[110]^x[85]^x[84]^x[74]^x[31]^x[20]^x[19]^x[8];
	y[19]=x[350]^x[339]^x[190]^x[184]^x[179]^x[178]^x[173]^x[172]^x[167]^x[161]^x[115]^x[109]^x[84]^x[83]^x[73]^x[30]^x[19]^x[18]^x[7];
	y[18]=x[349]^x[338]^x[189]^x[183]^x[178]^x[177]^x[172]^x[171]^x[166]^x[160]^x[114]^x[108]^x[83]^x[82]^x[72]^x[29]^x[18]^x[17]^x[6];
	y[17]=x[348]^x[337]^x[188]^x[182]^x[177]^x[176]^x[171]^x[165]^x[113]^x[107]^x[82]^x[81]^x[71]^x[28]^x[17]^x[16]^x[5];
	y[16]=x[347]^x[336]^x[187]^x[181]^x[176]^x[175]^x[170]^x[164]^x[112]^x[106]^x[81]^x[80]^x[70]^x[27]^x[16]^x[15]^x[4];
	y[15]=x[346]^x[335]^x[186]^x[180]^x[175]^x[174]^x[169]^x[163]^x[111]^x[105]^x[80]^x[79]^x[69]^x[26]^x[15]^x[14]^x[3];
	y[14]=x[345]^x[334]^x[185]^x[179]^x[174]^x[173]^x[168]^x[162]^x[110]^x[104]^x[79]^x[78]^x[68]^x[25]^x[14]^x[13]^x[2];
	y[13]=x[344]^x[333]^x[184]^x[178]^x[173]^x[172]^x[167]^x[161]^x[109]^x[103]^x[78]^x[77]^x[67]^x[24]^x[13]^x[12]^x[1];
	y[12]=x[343]^x[332]^x[183]^x[177]^x[172]^x[171]^x[166]^x[160]^x[108]^x[102]^x[77]^x[76]^x[66]^x[23]^x[12]^x[11]^x[0];
	y[11]=x[342]^x[331]^x[182]^x[176]^x[171]^x[165]^x[107]^x[101]^x[76]^x[75]^x[65]^x[22]^x[11];
	y[10]=x[341]^x[330]^x[181]^x[175]^x[170]^x[164]^x[106]^x[100]^x[75]^x[74]^x[64]^x[21]^x[10];
	y[9]=x[340]^x[329]^x[180]^x[174]^x[169]^x[163]^x[105]^x[99]^x[95]^x[73]^x[20]^x[9];
	y[8]=x[339]^x[328]^x[179]^x[173]^x[168]^x[162]^x[104]^x[98]^x[94]^x[72]^x[19]^x[8];
	y[7]=x[338]^x[327]^x[178]^x[172]^x[167]^x[161]^x[103]^x[97]^x[93]^x[71]^x[18]^x[7];
	y[6]=x[337]^x[326]^x[177]^x[171]^x[166]^x[160]^x[102]^x[96]^x[92]^x[70]^x[17]^x[6];
	y[5]=x[336]^x[325]^x[245]^x[234]^x[176]^x[165]^x[101]^x[91]^x[69]^x[16]^x[10]^x[5]^x[4];
	y[4]=x[335]^x[324]^x[244]^x[233]^x[175]^x[164]^x[100]^x[90]^x[68]^x[15]^x[9]^x[4]^x[3];
	y[3]=x[334]^x[323]^x[243]^x[232]^x[174]^x[163]^x[99]^x[89]^x[67]^x[14]^x[8]^x[3]^x[2];
	y[2]=x[333]^x[322]^x[242]^x[231]^x[173]^x[162]^x[98]^x[88]^x[66]^x[13]^x[7]^x[2]^x[1];
	y[1]=x[332]^x[321]^x[241]^x[230]^x[172]^x[161]^x[97]^x[87]^x[65]^x[12]^x[6]^x[1]^x[0];
	y[0]=x[331]^x[320]^x[240]^x[229]^x[171]^x[160]^x[96]^x[86]^x[64]^x[11]^x[5]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint22(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[373]^x[372]^x[371]^x[363]^x[361]^x[352]^x[319]^x[309]^x[306]^x[298]^x[295]^x[95]^x[89]^x[71]^x[65]^x[63]^x[53]^x[43]^x[32];
	y[30]=x[383]^x[382]^x[372]^x[371]^x[370]^x[360]^x[318]^x[308]^x[305]^x[297]^x[294]^x[94]^x[88]^x[70]^x[64]^x[63]^x[62]^x[52];
	y[29]=x[382]^x[381]^x[371]^x[370]^x[369]^x[359]^x[317]^x[307]^x[304]^x[296]^x[293]^x[93]^x[87]^x[69]^x[62]^x[61]^x[51];
	y[28]=x[381]^x[380]^x[370]^x[369]^x[368]^x[358]^x[316]^x[306]^x[303]^x[295]^x[292]^x[92]^x[86]^x[68]^x[61]^x[60]^x[50];
	y[27]=x[380]^x[379]^x[369]^x[368]^x[367]^x[357]^x[315]^x[305]^x[302]^x[294]^x[291]^x[91]^x[85]^x[67]^x[60]^x[59]^x[49];
	y[26]=x[383]^x[379]^x[378]^x[377]^x[368]^x[367]^x[366]^x[356]^x[314]^x[304]^x[301]^x[293]^x[290]^x[223]^x[147]^x[90]^x[84]^x[66]^x[59]^x[58]^x[48];
	y[25]=x[382]^x[378]^x[377]^x[376]^x[367]^x[366]^x[365]^x[355]^x[313]^x[303]^x[300]^x[292]^x[289]^x[222]^x[146]^x[89]^x[83]^x[65]^x[58]^x[57]^x[47];
	y[24]=x[381]^x[377]^x[376]^x[375]^x[366]^x[365]^x[364]^x[354]^x[312]^x[302]^x[299]^x[291]^x[288]^x[221]^x[145]^x[88]^x[82]^x[64]^x[57]^x[56]^x[46];
	y[23]=x[380]^x[376]^x[375]^x[374]^x[365]^x[364]^x[363]^x[353]^x[311]^x[301]^x[290]^x[220]^x[144]^x[87]^x[81]^x[56]^x[55]^x[45];
	y[22]=x[379]^x[375]^x[374]^x[373]^x[364]^x[363]^x[362]^x[352]^x[310]^x[300]^x[289]^x[219]^x[143]^x[86]^x[80]^x[55]^x[54]^x[44];
	y[21]=x[378]^x[374]^x[373]^x[372]^x[363]^x[361]^x[309]^x[299]^x[288]^x[218]^x[142]^x[85]^x[79]^x[54]^x[53]^x[43];
	y[20]=x[382]^x[373]^x[372]^x[362]^x[360]^x[319]^x[308]^x[84]^x[78]^x[53]^x[52]^x[42];
	y[19]=x[381]^x[372]^x[371]^x[361]^x[359]^x[318]^x[307]^x[83]^x[77]^x[52]^x[51]^x[41];
	y[18]=x[380]^x[371]^x[370]^x[360]^x[358]^x[317]^x[306]^x[82]^x[76]^x[51]^x[50]^x[40];
	y[17]=x[379]^x[370]^x[369]^x[359]^x[357]^x[316]^x[305]^x[138]^x[81]^x[75]^x[50]^x[49]^x[39];
	y[16]=x[378]^x[369]^x[368]^x[358]^x[356]^x[315]^x[304]^x[137]^x[80]^x[74]^x[49]^x[48]^x[38];
	y[15]=x[377]^x[368]^x[367]^x[357]^x[355]^x[314]^x[303]^x[136]^x[79]^x[73]^x[48]^x[47]^x[37];
	y[14]=x[376]^x[367]^x[366]^x[356]^x[354]^x[313]^x[302]^x[135]^x[78]^x[72]^x[47]^x[46]^x[36];
	y[13]=x[375]^x[366]^x[365]^x[355]^x[353]^x[312]^x[301]^x[134]^x[77]^x[71]^x[46]^x[45]^x[35];
	y[12]=x[374]^x[365]^x[364]^x[354]^x[352]^x[311]^x[300]^x[133]^x[76]^x[70]^x[45]^x[44]^x[34];
	y[11]=x[364]^x[363]^x[353]^x[310]^x[299]^x[75]^x[69]^x[44]^x[43]^x[33];
	y[10]=x[363]^x[362]^x[352]^x[309]^x[298]^x[74]^x[68]^x[43]^x[42]^x[32];
	y[9]=x[383]^x[361]^x[308]^x[297]^x[73]^x[67]^x[63]^x[41];
	y[8]=x[382]^x[360]^x[307]^x[296]^x[72]^x[66]^x[62]^x[40];
	y[7]=x[381]^x[359]^x[306]^x[295]^x[71]^x[65]^x[61]^x[39];
	y[6]=x[380]^x[358]^x[305]^x[294]^x[70]^x[64]^x[60]^x[38];
	y[5]=x[379]^x[373]^x[367]^x[362]^x[357]^x[356]^x[304]^x[293]^x[213]^x[202]^x[69]^x[59]^x[37];
	y[4]=x[378]^x[372]^x[366]^x[361]^x[356]^x[355]^x[303]^x[292]^x[212]^x[201]^x[68]^x[58]^x[36];
	y[3]=x[377]^x[371]^x[365]^x[360]^x[355]^x[354]^x[302]^x[291]^x[211]^x[200]^x[67]^x[57]^x[35];
	y[2]=x[376]^x[370]^x[364]^x[359]^x[354]^x[353]^x[301]^x[290]^x[210]^x[199]^x[66]^x[56]^x[34];
	y[1]=x[375]^x[369]^x[363]^x[358]^x[353]^x[352]^x[300]^x[289]^x[209]^x[198]^x[65]^x[55]^x[33];
	y[0]=x[374]^x[368]^x[357]^x[352]^x[299]^x[288]^x[208]^x[197]^x[64]^x[54]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint23(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[341]^x[340]^x[339]^x[331]^x[329]^x[320]^x[287]^x[277]^x[274]^x[266]^x[263]^x[63]^x[57]^x[39]^x[33]^x[31]^x[21]^x[11]^x[0];
	y[30]=x[351]^x[350]^x[340]^x[339]^x[338]^x[328]^x[286]^x[276]^x[273]^x[265]^x[262]^x[62]^x[56]^x[38]^x[32]^x[31]^x[30]^x[20];
	y[29]=x[350]^x[349]^x[339]^x[338]^x[337]^x[327]^x[285]^x[275]^x[272]^x[264]^x[261]^x[61]^x[55]^x[37]^x[30]^x[29]^x[19];
	y[28]=x[349]^x[348]^x[338]^x[337]^x[336]^x[326]^x[284]^x[274]^x[271]^x[263]^x[260]^x[60]^x[54]^x[36]^x[29]^x[28]^x[18];
	y[27]=x[348]^x[347]^x[337]^x[336]^x[335]^x[325]^x[283]^x[273]^x[270]^x[262]^x[259]^x[59]^x[53]^x[35]^x[28]^x[27]^x[17];
	y[26]=x[351]^x[347]^x[346]^x[345]^x[336]^x[335]^x[334]^x[324]^x[282]^x[272]^x[269]^x[261]^x[258]^x[191]^x[115]^x[58]^x[52]^x[34]^x[27]^x[26]^x[16];
	y[25]=x[350]^x[346]^x[345]^x[344]^x[335]^x[334]^x[333]^x[323]^x[281]^x[271]^x[268]^x[260]^x[257]^x[190]^x[114]^x[57]^x[51]^x[33]^x[26]^x[25]^x[15];
	y[24]=x[349]^x[345]^x[344]^x[343]^x[334]^x[333]^x[332]^x[322]^x[280]^x[270]^x[267]^x[259]^x[256]^x[189]^x[113]^x[56]^x[50]^x[32]^x[25]^x[24]^x[14];
	y[23]=x[348]^x[344]^x[343]^x[342]^x[333]^x[332]^x[331]^x[321]^x[279]^x[269]^x[258]^x[188]^x[112]^x[55]^x[49]^x[24]^x[23]^x[13];
	y[22]=x[347]^x[343]^x[342]^x[341]^x[332]^x[331]^x[330]^x[320]^x[278]^x[268]^x[257]^x[187]^x[111]^x[54]^x[48]^x[23]^x[22]^x[12];
	y[21]=x[346]^x[342]^x[341]^x[340]^x[331]^x[329]^x[277]^x[267]^x[256]^x[186]^x[110]^x[53]^x[47]^x[22]^x[21]^x[11];
	y[20]=x[350]^x[341]^x[340]^x[330]^x[328]^x[287]^x[276]^x[52]^x[46]^x[21]^x[20]^x[10];
	y[19]=x[349]^x[340]^x[339]^x[329]^x[327]^x[286]^x[275]^x[51]^x[45]^x[20]^x[19]^x[9];
	y[18]=x[348]^x[339]^x[338]^x[328]^x[326]^x[285]^x[274]^x[50]^x[44]^x[19]^x[18]^x[8];
	y[17]=x[347]^x[338]^x[337]^x[327]^x[325]^x[284]^x[273]^x[106]^x[49]^x[43]^x[18]^x[17]^x[7];
	y[16]=x[346]^x[337]^x[336]^x[326]^x[324]^x[283]^x[272]^x[105]^x[48]^x[42]^x[17]^x[16]^x[6];
	y[15]=x[345]^x[336]^x[335]^x[325]^x[323]^x[282]^x[271]^x[104]^x[47]^x[41]^x[16]^x[15]^x[5];
	y[14]=x[344]^x[335]^x[334]^x[324]^x[322]^x[281]^x[270]^x[103]^x[46]^x[40]^x[15]^x[14]^x[4];
	y[13]=x[343]^x[334]^x[333]^x[323]^x[321]^x[280]^x[269]^x[102]^x[45]^x[39]^x[14]^x[13]^x[3];
	y[12]=x[342]^x[333]^x[332]^x[322]^x[320]^x[279]^x[268]^x[101]^x[44]^x[38]^x[13]^x[12]^x[2];
	y[11]=x[332]^x[331]^x[321]^x[278]^x[267]^x[43]^x[37]^x[12]^x[11]^x[1];
	y[10]=x[331]^x[330]^x[320]^x[277]^x[266]^x[42]^x[36]^x[11]^x[10]^x[0];
	y[9]=x[351]^x[329]^x[276]^x[265]^x[41]^x[35]^x[31]^x[9];
	y[8]=x[350]^x[328]^x[275]^x[264]^x[40]^x[34]^x[30]^x[8];
	y[7]=x[349]^x[327]^x[274]^x[263]^x[39]^x[33]^x[29]^x[7];
	y[6]=x[348]^x[326]^x[273]^x[262]^x[38]^x[32]^x[28]^x[6];
	y[5]=x[347]^x[341]^x[335]^x[330]^x[325]^x[324]^x[272]^x[261]^x[181]^x[170]^x[37]^x[27]^x[5];
	y[4]=x[346]^x[340]^x[334]^x[329]^x[324]^x[323]^x[271]^x[260]^x[180]^x[169]^x[36]^x[26]^x[4];
	y[3]=x[345]^x[339]^x[333]^x[328]^x[323]^x[322]^x[270]^x[259]^x[179]^x[168]^x[35]^x[25]^x[3];
	y[2]=x[344]^x[338]^x[332]^x[327]^x[322]^x[321]^x[269]^x[258]^x[178]^x[167]^x[34]^x[24]^x[2];
	y[1]=x[343]^x[337]^x[331]^x[326]^x[321]^x[320]^x[268]^x[257]^x[177]^x[166]^x[33]^x[23]^x[1];
	y[0]=x[342]^x[336]^x[325]^x[320]^x[267]^x[256]^x[176]^x[165]^x[32]^x[22]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint24(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[374]^x[363]^x[362]^x[319]^x[309]^x[308]^x[307]^x[299]^x[297]^x[288]^x[255]^x[245]^x[242]^x[234]^x[231]^x[159]^x[153]^x[149]^x[143]^x[139]^x[133]^x[128]^x[31]^x[25]^x[7]^x[1];
	y[30]=x[382]^x[373]^x[362]^x[361]^x[319]^x[318]^x[308]^x[307]^x[306]^x[296]^x[254]^x[244]^x[241]^x[233]^x[230]^x[159]^x[158]^x[153]^x[152]^x[148]^x[142]^x[30]^x[24]^x[6]^x[0];
	y[29]=x[381]^x[372]^x[361]^x[360]^x[318]^x[317]^x[307]^x[306]^x[305]^x[295]^x[253]^x[243]^x[240]^x[232]^x[229]^x[158]^x[157]^x[152]^x[151]^x[147]^x[141]^x[29]^x[23]^x[5];
	y[28]=x[380]^x[371]^x[360]^x[359]^x[317]^x[316]^x[306]^x[305]^x[304]^x[294]^x[252]^x[242]^x[239]^x[231]^x[228]^x[157]^x[156]^x[151]^x[150]^x[146]^x[140]^x[28]^x[22]^x[4];
	y[27]=x[379]^x[370]^x[359]^x[358]^x[316]^x[315]^x[305]^x[304]^x[303]^x[293]^x[251]^x[241]^x[238]^x[230]^x[227]^x[156]^x[155]^x[150]^x[149]^x[145]^x[139]^x[27]^x[21]^x[3];
	y[26]=x[378]^x[369]^x[358]^x[357]^x[319]^x[315]^x[314]^x[313]^x[304]^x[303]^x[302]^x[292]^x[250]^x[240]^x[237]^x[229]^x[226]^x[159]^x[155]^x[154]^x[149]^x[148]^x[144]^x[138]^x[83]^x[26]^x[20]^x[2];
	y[25]=x[377]^x[368]^x[357]^x[356]^x[318]^x[314]^x[313]^x[312]^x[303]^x[302]^x[301]^x[291]^x[249]^x[239]^x[236]^x[228]^x[225]^x[158]^x[154]^x[153]^x[148]^x[147]^x[143]^x[137]^x[82]^x[25]^x[19]^x[1];
	y[24]=x[376]^x[367]^x[356]^x[355]^x[317]^x[313]^x[312]^x[311]^x[302]^x[301]^x[300]^x[290]^x[248]^x[238]^x[235]^x[227]^x[224]^x[157]^x[153]^x[152]^x[147]^x[146]^x[142]^x[136]^x[81]^x[24]^x[18]^x[0];
	y[23]=x[375]^x[366]^x[355]^x[354]^x[316]^x[312]^x[311]^x[310]^x[301]^x[300]^x[299]^x[289]^x[247]^x[237]^x[226]^x[156]^x[152]^x[151]^x[146]^x[145]^x[141]^x[135]^x[80]^x[23]^x[17];
	y[22]=x[374]^x[365]^x[354]^x[353]^x[315]^x[311]^x[310]^x[309]^x[300]^x[299]^x[298]^x[288]^x[246]^x[236]^x[225]^x[155]^x[151]^x[150]^x[145]^x[144]^x[140]^x[134]^x[79]^x[22]^x[16];
	y[21]=x[373]^x[364]^x[353]^x[352]^x[314]^x[310]^x[309]^x[308]^x[299]^x[297]^x[245]^x[235]^x[224]^x[154]^x[150]^x[149]^x[144]^x[143]^x[139]^x[133]^x[78]^x[21]^x[15];
	y[20]=x[383]^x[372]^x[363]^x[362]^x[352]^x[318]^x[309]^x[308]^x[298]^x[296]^x[255]^x[244]^x[149]^x[148]^x[143]^x[142]^x[138]^x[132]^x[20]^x[14];
	y[19]=x[383]^x[382]^x[371]^x[361]^x[317]^x[308]^x[307]^x[297]^x[295]^x[254]^x[243]^x[148]^x[147]^x[142]^x[141]^x[137]^x[131]^x[19]^x[13];
	y[18]=x[382]^x[381]^x[370]^x[360]^x[316]^x[307]^x[306]^x[296]^x[294]^x[253]^x[242]^x[147]^x[146]^x[141]^x[140]^x[136]^x[130]^x[18]^x[12];
	y[17]=x[381]^x[380]^x[369]^x[359]^x[315]^x[306]^x[305]^x[295]^x[293]^x[252]^x[241]^x[146]^x[145]^x[140]^x[139]^x[135]^x[129]^x[74]^x[17]^x[11];
	y[16]=x[380]^x[379]^x[368]^x[358]^x[314]^x[305]^x[304]^x[294]^x[292]^x[251]^x[240]^x[145]^x[144]^x[139]^x[138]^x[134]^x[128]^x[73]^x[16]^x[10];
	y[15]=x[379]^x[378]^x[367]^x[357]^x[313]^x[304]^x[303]^x[293]^x[291]^x[250]^x[239]^x[144]^x[143]^x[138]^x[137]^x[133]^x[72]^x[15]^x[9];
	y[14]=x[378]^x[377]^x[366]^x[356]^x[312]^x[303]^x[302]^x[292]^x[290]^x[249]^x[238]^x[143]^x[142]^x[137]^x[136]^x[132]^x[71]^x[14]^x[8];
	y[13]=x[377]^x[376]^x[365]^x[355]^x[311]^x[302]^x[301]^x[291]^x[289]^x[248]^x[237]^x[142]^x[141]^x[136]^x[135]^x[131]^x[70]^x[13]^x[7];
	y[12]=x[376]^x[375]^x[364]^x[354]^x[310]^x[301]^x[300]^x[290]^x[288]^x[247]^x[236]^x[141]^x[140]^x[135]^x[134]^x[130]^x[69]^x[12]^x[6];
	y[11]=x[375]^x[374]^x[363]^x[353]^x[300]^x[299]^x[289]^x[246]^x[235]^x[140]^x[139]^x[134]^x[133]^x[129]^x[11]^x[5];
	y[10]=x[374]^x[373]^x[362]^x[352]^x[299]^x[298]^x[288]^x[245]^x[234]^x[139]^x[138]^x[133]^x[132]^x[128]^x[10]^x[4];
	y[9]=x[383]^x[373]^x[372]^x[362]^x[361]^x[319]^x[297]^x[244]^x[233]^x[159]^x[153]^x[137]^x[131]^x[9]^x[3];
	y[8]=x[382]^x[372]^x[371]^x[361]^x[360]^x[318]^x[296]^x[243]^x[232]^x[158]^x[152]^x[136]^x[130]^x[8]^x[2];
	y[7]=x[381]^x[371]^x[370]^x[360]^x[359]^x[317]^x[295]^x[242]^x[231]^x[157]^x[151]^x[135]^x[129]^x[7]^x[1];
	y[6]=x[380]^x[370]^x[369]^x[359]^x[358]^x[316]^x[294]^x[241]^x[230]^x[156]^x[150]^x[134]^x[128]^x[6]^x[0];
	y[5]=x[379]^x[369]^x[368]^x[358]^x[357]^x[315]^x[309]^x[303]^x[298]^x[293]^x[292]^x[240]^x[229]^x[155]^x[138]^x[133]^x[5];
	y[4]=x[378]^x[368]^x[367]^x[357]^x[356]^x[314]^x[308]^x[302]^x[297]^x[292]^x[291]^x[239]^x[228]^x[154]^x[137]^x[132]^x[4];
	y[3]=x[377]^x[367]^x[366]^x[356]^x[355]^x[313]^x[307]^x[301]^x[296]^x[291]^x[290]^x[238]^x[227]^x[153]^x[136]^x[131]^x[3];
	y[2]=x[376]^x[366]^x[365]^x[355]^x[354]^x[312]^x[306]^x[300]^x[295]^x[290]^x[289]^x[237]^x[226]^x[152]^x[135]^x[130]^x[2];
	y[1]=x[375]^x[365]^x[364]^x[354]^x[353]^x[311]^x[305]^x[299]^x[294]^x[289]^x[288]^x[236]^x[225]^x[151]^x[134]^x[129]^x[1];
	y[0]=x[374]^x[364]^x[363]^x[353]^x[352]^x[310]^x[304]^x[293]^x[288]^x[235]^x[224]^x[150]^x[133]^x[128]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint25(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[377]^x[373]^x[370]^x[367]^x[364]^x[362]^x[359]^x[356]^x[353]^x[351]^x[342]^x[331]^x[330]^x[287]^x[277]^x[276]^x[275]^x[267]^x[265]^x[256]^x[223]^x[213]^x[210]^x[202]^x[199]^x[159]^x[147]^x[135]^x[127]^x[121]^x[117]^x[111]^x[107]^x[101]^x[96];
	y[30]=x[382]^x[376]^x[372]^x[369]^x[366]^x[363]^x[361]^x[358]^x[355]^x[352]^x[350]^x[341]^x[330]^x[329]^x[287]^x[286]^x[276]^x[275]^x[274]^x[264]^x[222]^x[212]^x[209]^x[201]^x[198]^x[158]^x[146]^x[134]^x[127]^x[126]^x[121]^x[120]^x[116]^x[110];
	y[29]=x[381]^x[375]^x[371]^x[368]^x[365]^x[360]^x[357]^x[354]^x[349]^x[340]^x[329]^x[328]^x[286]^x[285]^x[275]^x[274]^x[273]^x[263]^x[221]^x[211]^x[208]^x[200]^x[197]^x[157]^x[145]^x[133]^x[126]^x[125]^x[120]^x[119]^x[115]^x[109];
	y[28]=x[380]^x[374]^x[370]^x[367]^x[364]^x[359]^x[356]^x[353]^x[348]^x[339]^x[328]^x[327]^x[285]^x[284]^x[274]^x[273]^x[272]^x[262]^x[220]^x[210]^x[207]^x[199]^x[196]^x[156]^x[144]^x[132]^x[125]^x[124]^x[119]^x[118]^x[114]^x[108];
	y[27]=x[379]^x[373]^x[369]^x[366]^x[363]^x[358]^x[355]^x[352]^x[347]^x[338]^x[327]^x[326]^x[284]^x[283]^x[273]^x[272]^x[271]^x[261]^x[219]^x[209]^x[206]^x[198]^x[195]^x[155]^x[143]^x[131]^x[124]^x[123]^x[118]^x[117]^x[113]^x[107];
	y[26]=x[383]^x[378]^x[372]^x[368]^x[365]^x[357]^x[354]^x[346]^x[337]^x[326]^x[325]^x[287]^x[283]^x[282]^x[281]^x[272]^x[271]^x[270]^x[260]^x[218]^x[208]^x[205]^x[197]^x[194]^x[154]^x[142]^x[130]^x[127]^x[123]^x[122]^x[117]^x[116]^x[112]^x[106]^x[51];
	y[25]=x[382]^x[377]^x[371]^x[367]^x[364]^x[356]^x[353]^x[345]^x[336]^x[325]^x[324]^x[286]^x[282]^x[281]^x[280]^x[271]^x[270]^x[269]^x[259]^x[217]^x[207]^x[204]^x[196]^x[193]^x[153]^x[141]^x[129]^x[126]^x[122]^x[121]^x[116]^x[115]^x[111]^x[105]^x[50];
	y[24]=x[381]^x[376]^x[370]^x[366]^x[363]^x[355]^x[352]^x[344]^x[335]^x[324]^x[323]^x[285]^x[281]^x[280]^x[279]^x[270]^x[269]^x[268]^x[258]^x[216]^x[206]^x[203]^x[195]^x[192]^x[152]^x[140]^x[128]^x[125]^x[121]^x[120]^x[115]^x[114]^x[110]^x[104]^x[49];
	y[23]=x[380]^x[375]^x[369]^x[365]^x[354]^x[343]^x[334]^x[323]^x[322]^x[284]^x[280]^x[279]^x[278]^x[269]^x[268]^x[267]^x[257]^x[215]^x[205]^x[194]^x[151]^x[139]^x[124]^x[120]^x[119]^x[114]^x[113]^x[109]^x[103]^x[48];
	y[22]=x[379]^x[374]^x[368]^x[364]^x[353]^x[342]^x[333]^x[322]^x[321]^x[283]^x[279]^x[278]^x[277]^x[268]^x[267]^x[266]^x[256]^x[214]^x[204]^x[193]^x[150]^x[138]^x[123]^x[119]^x[118]^x[113]^x[112]^x[108]^x[102]^x[47];
	y[21]=x[378]^x[373]^x[367]^x[363]^x[352]^x[341]^x[332]^x[321]^x[320]^x[282]^x[278]^x[277]^x[276]^x[267]^x[265]^x[213]^x[203]^x[192]^x[149]^x[137]^x[122]^x[118]^x[117]^x[112]^x[111]^x[107]^x[101]^x[46];
	y[20]=x[383]^x[377]^x[372]^x[366]^x[351]^x[340]^x[331]^x[330]^x[320]^x[286]^x[277]^x[276]^x[266]^x[264]^x[223]^x[212]^x[148]^x[136]^x[117]^x[116]^x[111]^x[110]^x[106]^x[100];
	y[19]=x[382]^x[376]^x[371]^x[365]^x[351]^x[350]^x[339]^x[329]^x[285]^x[276]^x[275]^x[265]^x[263]^x[222]^x[211]^x[147]^x[135]^x[116]^x[115]^x[110]^x[109]^x[105]^x[99];
	y[18]=x[381]^x[375]^x[370]^x[364]^x[350]^x[349]^x[338]^x[328]^x[284]^x[275]^x[274]^x[264]^x[262]^x[221]^x[210]^x[146]^x[134]^x[115]^x[114]^x[109]^x[108]^x[104]^x[98];
	y[17]=x[380]^x[374]^x[369]^x[363]^x[349]^x[348]^x[337]^x[327]^x[283]^x[274]^x[273]^x[263]^x[261]^x[220]^x[209]^x[145]^x[133]^x[114]^x[113]^x[108]^x[107]^x[103]^x[97]^x[42];
	y[16]=x[379]^x[373]^x[368]^x[362]^x[348]^x[347]^x[336]^x[326]^x[282]^x[273]^x[272]^x[262]^x[260]^x[219]^x[208]^x[144]^x[132]^x[113]^x[112]^x[107]^x[106]^x[102]^x[96]^x[41];
	y[15]=x[378]^x[372]^x[367]^x[361]^x[347]^x[346]^x[335]^x[325]^x[281]^x[272]^x[271]^x[261]^x[259]^x[218]^x[207]^x[143]^x[131]^x[112]^x[111]^x[106]^x[105]^x[101]^x[40];
	y[14]=x[377]^x[371]^x[366]^x[360]^x[346]^x[345]^x[334]^x[324]^x[280]^x[271]^x[270]^x[260]^x[258]^x[217]^x[206]^x[142]^x[130]^x[111]^x[110]^x[105]^x[104]^x[100]^x[39];
	y[13]=x[376]^x[370]^x[365]^x[359]^x[345]^x[344]^x[333]^x[323]^x[279]^x[270]^x[269]^x[259]^x[257]^x[216]^x[205]^x[141]^x[129]^x[110]^x[109]^x[104]^x[103]^x[99]^x[38];
	y[12]=x[375]^x[369]^x[364]^x[358]^x[344]^x[343]^x[332]^x[322]^x[278]^x[269]^x[268]^x[258]^x[256]^x[215]^x[204]^x[140]^x[128]^x[109]^x[108]^x[103]^x[102]^x[98]^x[37];
	y[11]=x[374]^x[368]^x[363]^x[357]^x[343]^x[342]^x[331]^x[321]^x[268]^x[267]^x[257]^x[214]^x[203]^x[139]^x[108]^x[107]^x[102]^x[101]^x[97];
	y[10]=x[373]^x[367]^x[362]^x[356]^x[342]^x[341]^x[330]^x[320]^x[267]^x[266]^x[256]^x[213]^x[202]^x[138]^x[107]^x[106]^x[101]^x[100]^x[96];
	y[9]=x[372]^x[366]^x[361]^x[355]^x[351]^x[341]^x[340]^x[330]^x[329]^x[287]^x[265]^x[212]^x[201]^x[137]^x[127]^x[121]^x[105]^x[99];
	y[8]=x[371]^x[365]^x[360]^x[354]^x[350]^x[340]^x[339]^x[329]^x[328]^x[286]^x[264]^x[211]^x[200]^x[136]^x[126]^x[120]^x[104]^x[98];
	y[7]=x[370]^x[364]^x[359]^x[353]^x[349]^x[339]^x[338]^x[328]^x[327]^x[285]^x[263]^x[210]^x[199]^x[135]^x[125]^x[119]^x[103]^x[97];
	y[6]=x[369]^x[363]^x[358]^x[352]^x[348]^x[338]^x[337]^x[327]^x[326]^x[284]^x[262]^x[209]^x[198]^x[134]^x[124]^x[118]^x[102]^x[96];
	y[5]=x[368]^x[357]^x[347]^x[337]^x[336]^x[326]^x[325]^x[283]^x[277]^x[271]^x[266]^x[261]^x[260]^x[208]^x[197]^x[133]^x[123]^x[106]^x[101];
	y[4]=x[367]^x[356]^x[346]^x[336]^x[335]^x[325]^x[324]^x[282]^x[276]^x[270]^x[265]^x[260]^x[259]^x[207]^x[196]^x[132]^x[122]^x[105]^x[100];
	y[3]=x[366]^x[355]^x[345]^x[335]^x[334]^x[324]^x[323]^x[281]^x[275]^x[269]^x[264]^x[259]^x[258]^x[206]^x[195]^x[131]^x[121]^x[104]^x[99];
	y[2]=x[365]^x[354]^x[344]^x[334]^x[333]^x[323]^x[322]^x[280]^x[274]^x[268]^x[263]^x[258]^x[257]^x[205]^x[194]^x[130]^x[120]^x[103]^x[98];
	y[1]=x[364]^x[353]^x[343]^x[333]^x[332]^x[322]^x[321]^x[279]^x[273]^x[267]^x[262]^x[257]^x[256]^x[204]^x[193]^x[129]^x[119]^x[102]^x[97];
	y[0]=x[363]^x[352]^x[342]^x[332]^x[331]^x[321]^x[320]^x[278]^x[272]^x[261]^x[256]^x[203]^x[192]^x[128]^x[118]^x[101]^x[96];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint26(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[345]^x[341]^x[338]^x[335]^x[332]^x[330]^x[327]^x[324]^x[321]^x[319]^x[310]^x[299]^x[298]^x[255]^x[245]^x[244]^x[243]^x[235]^x[233]^x[224]^x[191]^x[181]^x[178]^x[170]^x[167]^x[127]^x[115]^x[103]^x[95]^x[89]^x[85]^x[79]^x[75]^x[69]^x[64];
	y[30]=x[350]^x[344]^x[340]^x[337]^x[334]^x[331]^x[329]^x[326]^x[323]^x[320]^x[318]^x[309]^x[298]^x[297]^x[255]^x[254]^x[244]^x[243]^x[242]^x[232]^x[190]^x[180]^x[177]^x[169]^x[166]^x[126]^x[114]^x[102]^x[95]^x[94]^x[89]^x[88]^x[84]^x[78];
	y[29]=x[349]^x[343]^x[339]^x[336]^x[333]^x[328]^x[325]^x[322]^x[317]^x[308]^x[297]^x[296]^x[254]^x[253]^x[243]^x[242]^x[241]^x[231]^x[189]^x[179]^x[176]^x[168]^x[165]^x[125]^x[113]^x[101]^x[94]^x[93]^x[88]^x[87]^x[83]^x[77];
	y[28]=x[348]^x[342]^x[338]^x[335]^x[332]^x[327]^x[324]^x[321]^x[316]^x[307]^x[296]^x[295]^x[253]^x[252]^x[242]^x[241]^x[240]^x[230]^x[188]^x[178]^x[175]^x[167]^x[164]^x[124]^x[112]^x[100]^x[93]^x[92]^x[87]^x[86]^x[82]^x[76];
	y[27]=x[347]^x[341]^x[337]^x[334]^x[331]^x[326]^x[323]^x[320]^x[315]^x[306]^x[295]^x[294]^x[252]^x[251]^x[241]^x[240]^x[239]^x[229]^x[187]^x[177]^x[174]^x[166]^x[163]^x[123]^x[111]^x[99]^x[92]^x[91]^x[86]^x[85]^x[81]^x[75];
	y[26]=x[351]^x[346]^x[340]^x[336]^x[333]^x[325]^x[322]^x[314]^x[305]^x[294]^x[293]^x[255]^x[251]^x[250]^x[249]^x[240]^x[239]^x[238]^x[228]^x[186]^x[176]^x[173]^x[165]^x[162]^x[122]^x[110]^x[98]^x[95]^x[91]^x[90]^x[85]^x[84]^x[80]^x[74]^x[19];
	y[25]=x[350]^x[345]^x[339]^x[335]^x[332]^x[324]^x[321]^x[313]^x[304]^x[293]^x[292]^x[254]^x[250]^x[249]^x[248]^x[239]^x[238]^x[237]^x[227]^x[185]^x[175]^x[172]^x[164]^x[161]^x[121]^x[109]^x[97]^x[94]^x[90]^x[89]^x[84]^x[83]^x[79]^x[73]^x[18];
	y[24]=x[349]^x[344]^x[338]^x[334]^x[331]^x[323]^x[320]^x[312]^x[303]^x[292]^x[291]^x[253]^x[249]^x[248]^x[247]^x[238]^x[237]^x[236]^x[226]^x[184]^x[174]^x[171]^x[163]^x[160]^x[120]^x[108]^x[96]^x[93]^x[89]^x[88]^x[83]^x[82]^x[78]^x[72]^x[17];
	y[23]=x[348]^x[343]^x[337]^x[333]^x[322]^x[311]^x[302]^x[291]^x[290]^x[252]^x[248]^x[247]^x[246]^x[237]^x[236]^x[235]^x[225]^x[183]^x[173]^x[162]^x[119]^x[107]^x[92]^x[88]^x[87]^x[82]^x[81]^x[77]^x[71]^x[16];
	y[22]=x[347]^x[342]^x[336]^x[332]^x[321]^x[310]^x[301]^x[290]^x[289]^x[251]^x[247]^x[246]^x[245]^x[236]^x[235]^x[234]^x[224]^x[182]^x[172]^x[161]^x[118]^x[106]^x[91]^x[87]^x[86]^x[81]^x[80]^x[76]^x[70]^x[15];
	y[21]=x[346]^x[341]^x[335]^x[331]^x[320]^x[309]^x[300]^x[289]^x[288]^x[250]^x[246]^x[245]^x[244]^x[235]^x[233]^x[181]^x[171]^x[160]^x[117]^x[105]^x[90]^x[86]^x[85]^x[80]^x[79]^x[75]^x[69]^x[14];
	y[20]=x[351]^x[345]^x[340]^x[334]^x[319]^x[308]^x[299]^x[298]^x[288]^x[254]^x[245]^x[244]^x[234]^x[232]^x[191]^x[180]^x[116]^x[104]^x[85]^x[84]^x[79]^x[78]^x[74]^x[68];
	y[19]=x[350]^x[344]^x[339]^x[333]^x[319]^x[318]^x[307]^x[297]^x[253]^x[244]^x[243]^x[233]^x[231]^x[190]^x[179]^x[115]^x[103]^x[84]^x[83]^x[78]^x[77]^x[73]^x[67];
	y[18]=x[349]^x[343]^x[338]^x[332]^x[318]^x[317]^x[306]^x[296]^x[252]^x[243]^x[242]^x[232]^x[230]^x[189]^x[178]^x[114]^x[102]^x[83]^x[82]^x[77]^x[76]^x[72]^x[66];
	y[17]=x[348]^x[342]^x[337]^x[331]^x[317]^x[316]^x[305]^x[295]^x[251]^x[242]^x[241]^x[231]^x[229]^x[188]^x[177]^x[113]^x[101]^x[82]^x[81]^x[76]^x[75]^x[71]^x[65]^x[10];
	y[16]=x[347]^x[341]^x[336]^x[330]^x[316]^x[315]^x[304]^x[294]^x[250]^x[241]^x[240]^x[230]^x[228]^x[187]^x[176]^x[112]^x[100]^x[81]^x[80]^x[75]^x[74]^x[70]^x[64]^x[9];
	y[15]=x[346]^x[340]^x[335]^x[329]^x[315]^x[314]^x[303]^x[293]^x[249]^x[240]^x[239]^x[229]^x[227]^x[186]^x[175]^x[111]^x[99]^x[80]^x[79]^x[74]^x[73]^x[69]^x[8];
	y[14]=x[345]^x[339]^x[334]^x[328]^x[314]^x[313]^x[302]^x[292]^x[248]^x[239]^x[238]^x[228]^x[226]^x[185]^x[174]^x[110]^x[98]^x[79]^x[78]^x[73]^x[72]^x[68]^x[7];
	y[13]=x[344]^x[338]^x[333]^x[327]^x[313]^x[312]^x[301]^x[291]^x[247]^x[238]^x[237]^x[227]^x[225]^x[184]^x[173]^x[109]^x[97]^x[78]^x[77]^x[72]^x[71]^x[67]^x[6];
	y[12]=x[343]^x[337]^x[332]^x[326]^x[312]^x[311]^x[300]^x[290]^x[246]^x[237]^x[236]^x[226]^x[224]^x[183]^x[172]^x[108]^x[96]^x[77]^x[76]^x[71]^x[70]^x[66]^x[5];
	y[11]=x[342]^x[336]^x[331]^x[325]^x[311]^x[310]^x[299]^x[289]^x[236]^x[235]^x[225]^x[182]^x[171]^x[107]^x[76]^x[75]^x[70]^x[69]^x[65];
	y[10]=x[341]^x[335]^x[330]^x[324]^x[310]^x[309]^x[298]^x[288]^x[235]^x[234]^x[224]^x[181]^x[170]^x[106]^x[75]^x[74]^x[69]^x[68]^x[64];
	y[9]=x[340]^x[334]^x[329]^x[323]^x[319]^x[309]^x[308]^x[298]^x[297]^x[255]^x[233]^x[180]^x[169]^x[105]^x[95]^x[89]^x[73]^x[67];
	y[8]=x[339]^x[333]^x[328]^x[322]^x[318]^x[308]^x[307]^x[297]^x[296]^x[254]^x[232]^x[179]^x[168]^x[104]^x[94]^x[88]^x[72]^x[66];
	y[7]=x[338]^x[332]^x[327]^x[321]^x[317]^x[307]^x[306]^x[296]^x[295]^x[253]^x[231]^x[178]^x[167]^x[103]^x[93]^x[87]^x[71]^x[65];
	y[6]=x[337]^x[331]^x[326]^x[320]^x[316]^x[306]^x[305]^x[295]^x[294]^x[252]^x[230]^x[177]^x[166]^x[102]^x[92]^x[86]^x[70]^x[64];
	y[5]=x[336]^x[325]^x[315]^x[305]^x[304]^x[294]^x[293]^x[251]^x[245]^x[239]^x[234]^x[229]^x[228]^x[176]^x[165]^x[101]^x[91]^x[74]^x[69];
	y[4]=x[335]^x[324]^x[314]^x[304]^x[303]^x[293]^x[292]^x[250]^x[244]^x[238]^x[233]^x[228]^x[227]^x[175]^x[164]^x[100]^x[90]^x[73]^x[68];
	y[3]=x[334]^x[323]^x[313]^x[303]^x[302]^x[292]^x[291]^x[249]^x[243]^x[237]^x[232]^x[227]^x[226]^x[174]^x[163]^x[99]^x[89]^x[72]^x[67];
	y[2]=x[333]^x[322]^x[312]^x[302]^x[301]^x[291]^x[290]^x[248]^x[242]^x[236]^x[231]^x[226]^x[225]^x[173]^x[162]^x[98]^x[88]^x[71]^x[66];
	y[1]=x[332]^x[321]^x[311]^x[301]^x[300]^x[290]^x[289]^x[247]^x[241]^x[235]^x[230]^x[225]^x[224]^x[172]^x[161]^x[97]^x[87]^x[70]^x[65];
	y[0]=x[331]^x[320]^x[310]^x[300]^x[299]^x[289]^x[288]^x[246]^x[240]^x[229]^x[224]^x[171]^x[160]^x[96]^x[86]^x[69]^x[64];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint27(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[319]^x[313]^x[309]^x[306]^x[303]^x[300]^x[298]^x[295]^x[292]^x[289]^x[287]^x[278]^x[267]^x[266]^x[223]^x[213]^x[212]^x[211]^x[203]^x[201]^x[192]^x[159]^x[149]^x[146]^x[138]^x[135]^x[95]^x[83]^x[71]^x[63]^x[57]^x[53]^x[47]^x[43]^x[37]^x[32];
	y[30]=x[318]^x[312]^x[308]^x[305]^x[302]^x[299]^x[297]^x[294]^x[291]^x[288]^x[286]^x[277]^x[266]^x[265]^x[223]^x[222]^x[212]^x[211]^x[210]^x[200]^x[158]^x[148]^x[145]^x[137]^x[134]^x[94]^x[82]^x[70]^x[63]^x[62]^x[57]^x[56]^x[52]^x[46];
	y[29]=x[317]^x[311]^x[307]^x[304]^x[301]^x[296]^x[293]^x[290]^x[285]^x[276]^x[265]^x[264]^x[222]^x[221]^x[211]^x[210]^x[209]^x[199]^x[157]^x[147]^x[144]^x[136]^x[133]^x[93]^x[81]^x[69]^x[62]^x[61]^x[56]^x[55]^x[51]^x[45];
	y[28]=x[316]^x[310]^x[306]^x[303]^x[300]^x[295]^x[292]^x[289]^x[284]^x[275]^x[264]^x[263]^x[221]^x[220]^x[210]^x[209]^x[208]^x[198]^x[156]^x[146]^x[143]^x[135]^x[132]^x[92]^x[80]^x[68]^x[61]^x[60]^x[55]^x[54]^x[50]^x[44];
	y[27]=x[315]^x[309]^x[305]^x[302]^x[299]^x[294]^x[291]^x[288]^x[283]^x[274]^x[263]^x[262]^x[220]^x[219]^x[209]^x[208]^x[207]^x[197]^x[155]^x[145]^x[142]^x[134]^x[131]^x[91]^x[79]^x[67]^x[60]^x[59]^x[54]^x[53]^x[49]^x[43];
	y[26]=x[382]^x[371]^x[319]^x[314]^x[308]^x[304]^x[301]^x[293]^x[290]^x[282]^x[273]^x[262]^x[261]^x[223]^x[219]^x[218]^x[217]^x[208]^x[207]^x[206]^x[196]^x[154]^x[147]^x[144]^x[133]^x[130]^x[90]^x[78]^x[66]^x[63]^x[59]^x[58]^x[53]^x[52]^x[48]^x[42];
	y[25]=x[381]^x[370]^x[318]^x[313]^x[307]^x[303]^x[300]^x[292]^x[289]^x[281]^x[272]^x[261]^x[260]^x[222]^x[218]^x[217]^x[216]^x[207]^x[206]^x[205]^x[195]^x[153]^x[146]^x[143]^x[132]^x[129]^x[89]^x[77]^x[65]^x[62]^x[58]^x[57]^x[52]^x[51]^x[47]^x[41];
	y[24]=x[380]^x[369]^x[317]^x[312]^x[306]^x[302]^x[299]^x[291]^x[288]^x[280]^x[271]^x[260]^x[259]^x[221]^x[217]^x[216]^x[215]^x[206]^x[205]^x[204]^x[194]^x[152]^x[145]^x[142]^x[131]^x[128]^x[88]^x[76]^x[64]^x[61]^x[57]^x[56]^x[51]^x[50]^x[46]^x[40];
	y[23]=x[379]^x[368]^x[316]^x[311]^x[305]^x[301]^x[290]^x[279]^x[270]^x[259]^x[258]^x[220]^x[216]^x[215]^x[214]^x[205]^x[204]^x[203]^x[193]^x[151]^x[144]^x[141]^x[138]^x[130]^x[87]^x[75]^x[60]^x[56]^x[55]^x[50]^x[49]^x[45]^x[39];
	y[22]=x[378]^x[367]^x[315]^x[310]^x[304]^x[300]^x[289]^x[278]^x[269]^x[258]^x[257]^x[219]^x[215]^x[214]^x[213]^x[204]^x[203]^x[202]^x[192]^x[150]^x[143]^x[140]^x[137]^x[129]^x[86]^x[74]^x[59]^x[55]^x[54]^x[49]^x[48]^x[44]^x[38];
	y[21]=x[377]^x[366]^x[314]^x[309]^x[303]^x[299]^x[288]^x[277]^x[268]^x[257]^x[256]^x[218]^x[214]^x[213]^x[212]^x[203]^x[201]^x[149]^x[142]^x[139]^x[136]^x[128]^x[85]^x[73]^x[58]^x[54]^x[53]^x[48]^x[47]^x[43]^x[37];
	y[20]=x[319]^x[313]^x[308]^x[302]^x[287]^x[276]^x[267]^x[266]^x[256]^x[222]^x[213]^x[212]^x[202]^x[200]^x[159]^x[148]^x[84]^x[72]^x[53]^x[52]^x[47]^x[46]^x[42]^x[36];
	y[19]=x[318]^x[312]^x[307]^x[301]^x[287]^x[286]^x[275]^x[265]^x[221]^x[212]^x[211]^x[201]^x[199]^x[158]^x[147]^x[83]^x[71]^x[52]^x[51]^x[46]^x[45]^x[41]^x[35];
	y[18]=x[317]^x[311]^x[306]^x[300]^x[286]^x[285]^x[274]^x[264]^x[220]^x[211]^x[210]^x[200]^x[198]^x[157]^x[146]^x[82]^x[70]^x[51]^x[50]^x[45]^x[44]^x[40]^x[34];
	y[17]=x[373]^x[362]^x[316]^x[310]^x[305]^x[299]^x[285]^x[284]^x[273]^x[263]^x[219]^x[210]^x[209]^x[199]^x[197]^x[156]^x[145]^x[138]^x[132]^x[81]^x[69]^x[50]^x[49]^x[44]^x[43]^x[39]^x[33];
	y[16]=x[372]^x[361]^x[315]^x[309]^x[304]^x[298]^x[284]^x[283]^x[272]^x[262]^x[218]^x[209]^x[208]^x[198]^x[196]^x[155]^x[144]^x[137]^x[131]^x[80]^x[68]^x[49]^x[48]^x[43]^x[42]^x[38]^x[32];
	y[15]=x[371]^x[360]^x[314]^x[308]^x[303]^x[297]^x[283]^x[282]^x[271]^x[261]^x[217]^x[208]^x[207]^x[197]^x[195]^x[154]^x[143]^x[136]^x[130]^x[79]^x[67]^x[48]^x[47]^x[42]^x[41]^x[37];
	y[14]=x[370]^x[359]^x[313]^x[307]^x[302]^x[296]^x[282]^x[281]^x[270]^x[260]^x[216]^x[207]^x[206]^x[196]^x[194]^x[153]^x[142]^x[135]^x[129]^x[78]^x[66]^x[47]^x[46]^x[41]^x[40]^x[36];
	y[13]=x[369]^x[358]^x[312]^x[306]^x[301]^x[295]^x[281]^x[280]^x[269]^x[259]^x[215]^x[206]^x[205]^x[195]^x[193]^x[152]^x[141]^x[134]^x[128]^x[77]^x[65]^x[46]^x[45]^x[40]^x[39]^x[35];
	y[12]=x[368]^x[357]^x[311]^x[305]^x[300]^x[294]^x[280]^x[279]^x[268]^x[258]^x[214]^x[205]^x[204]^x[194]^x[192]^x[151]^x[140]^x[133]^x[76]^x[64]^x[45]^x[44]^x[39]^x[38]^x[34];
	y[11]=x[310]^x[304]^x[299]^x[293]^x[279]^x[278]^x[267]^x[257]^x[204]^x[203]^x[193]^x[150]^x[139]^x[75]^x[44]^x[43]^x[38]^x[37]^x[33];
	y[10]=x[309]^x[303]^x[298]^x[292]^x[278]^x[277]^x[266]^x[256]^x[203]^x[202]^x[192]^x[149]^x[138]^x[74]^x[43]^x[42]^x[37]^x[36]^x[32];
	y[9]=x[308]^x[302]^x[297]^x[291]^x[287]^x[277]^x[276]^x[266]^x[265]^x[223]^x[201]^x[148]^x[137]^x[73]^x[63]^x[57]^x[41]^x[35];
	y[8]=x[307]^x[301]^x[296]^x[290]^x[286]^x[276]^x[275]^x[265]^x[264]^x[222]^x[200]^x[147]^x[136]^x[72]^x[62]^x[56]^x[40]^x[34];
	y[7]=x[306]^x[300]^x[295]^x[289]^x[285]^x[275]^x[274]^x[264]^x[263]^x[221]^x[199]^x[146]^x[135]^x[71]^x[61]^x[55]^x[39]^x[33];
	y[6]=x[305]^x[299]^x[294]^x[288]^x[284]^x[274]^x[273]^x[263]^x[262]^x[220]^x[198]^x[145]^x[134]^x[70]^x[60]^x[54]^x[38]^x[32];
	y[5]=x[304]^x[293]^x[283]^x[273]^x[272]^x[262]^x[261]^x[219]^x[213]^x[207]^x[202]^x[197]^x[196]^x[144]^x[133]^x[69]^x[59]^x[42]^x[37];
	y[4]=x[303]^x[292]^x[282]^x[272]^x[271]^x[261]^x[260]^x[218]^x[212]^x[206]^x[201]^x[196]^x[195]^x[143]^x[132]^x[68]^x[58]^x[41]^x[36];
	y[3]=x[302]^x[291]^x[281]^x[271]^x[270]^x[260]^x[259]^x[217]^x[211]^x[205]^x[200]^x[195]^x[194]^x[142]^x[131]^x[67]^x[57]^x[40]^x[35];
	y[2]=x[301]^x[290]^x[280]^x[270]^x[269]^x[259]^x[258]^x[216]^x[210]^x[204]^x[199]^x[194]^x[193]^x[141]^x[130]^x[66]^x[56]^x[39]^x[34];
	y[1]=x[300]^x[289]^x[279]^x[269]^x[268]^x[258]^x[257]^x[215]^x[209]^x[203]^x[198]^x[193]^x[192]^x[140]^x[129]^x[65]^x[55]^x[38]^x[33];
	y[0]=x[299]^x[288]^x[278]^x[268]^x[267]^x[257]^x[256]^x[214]^x[208]^x[197]^x[192]^x[139]^x[128]^x[64]^x[54]^x[37]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint28(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[287]^x[281]^x[277]^x[274]^x[271]^x[268]^x[266]^x[263]^x[260]^x[257]^x[255]^x[246]^x[235]^x[234]^x[191]^x[181]^x[180]^x[179]^x[171]^x[169]^x[160]^x[127]^x[117]^x[114]^x[106]^x[103]^x[63]^x[51]^x[39]^x[31]^x[25]^x[21]^x[15]^x[11]^x[5]^x[0];
	y[30]=x[286]^x[280]^x[276]^x[273]^x[270]^x[267]^x[265]^x[262]^x[259]^x[256]^x[254]^x[245]^x[234]^x[233]^x[191]^x[190]^x[180]^x[179]^x[178]^x[168]^x[126]^x[116]^x[113]^x[105]^x[102]^x[62]^x[50]^x[38]^x[31]^x[30]^x[25]^x[24]^x[20]^x[14];
	y[29]=x[285]^x[279]^x[275]^x[272]^x[269]^x[264]^x[261]^x[258]^x[253]^x[244]^x[233]^x[232]^x[190]^x[189]^x[179]^x[178]^x[177]^x[167]^x[125]^x[115]^x[112]^x[104]^x[101]^x[61]^x[49]^x[37]^x[30]^x[29]^x[24]^x[23]^x[19]^x[13];
	y[28]=x[284]^x[278]^x[274]^x[271]^x[268]^x[263]^x[260]^x[257]^x[252]^x[243]^x[232]^x[231]^x[189]^x[188]^x[178]^x[177]^x[176]^x[166]^x[124]^x[114]^x[111]^x[103]^x[100]^x[60]^x[48]^x[36]^x[29]^x[28]^x[23]^x[22]^x[18]^x[12];
	y[27]=x[283]^x[277]^x[273]^x[270]^x[267]^x[262]^x[259]^x[256]^x[251]^x[242]^x[231]^x[230]^x[188]^x[187]^x[177]^x[176]^x[175]^x[165]^x[123]^x[113]^x[110]^x[102]^x[99]^x[59]^x[47]^x[35]^x[28]^x[27]^x[22]^x[21]^x[17]^x[11];
	y[26]=x[350]^x[339]^x[287]^x[282]^x[276]^x[272]^x[269]^x[261]^x[258]^x[250]^x[241]^x[230]^x[229]^x[191]^x[187]^x[186]^x[185]^x[176]^x[175]^x[174]^x[164]^x[122]^x[115]^x[112]^x[101]^x[98]^x[58]^x[46]^x[34]^x[31]^x[27]^x[26]^x[21]^x[20]^x[16]^x[10];
	y[25]=x[349]^x[338]^x[286]^x[281]^x[275]^x[271]^x[268]^x[260]^x[257]^x[249]^x[240]^x[229]^x[228]^x[190]^x[186]^x[185]^x[184]^x[175]^x[174]^x[173]^x[163]^x[121]^x[114]^x[111]^x[100]^x[97]^x[57]^x[45]^x[33]^x[30]^x[26]^x[25]^x[20]^x[19]^x[15]^x[9];
	y[24]=x[348]^x[337]^x[285]^x[280]^x[274]^x[270]^x[267]^x[259]^x[256]^x[248]^x[239]^x[228]^x[227]^x[189]^x[185]^x[184]^x[183]^x[174]^x[173]^x[172]^x[162]^x[120]^x[113]^x[110]^x[99]^x[96]^x[56]^x[44]^x[32]^x[29]^x[25]^x[24]^x[19]^x[18]^x[14]^x[8];
	y[23]=x[347]^x[336]^x[284]^x[279]^x[273]^x[269]^x[258]^x[247]^x[238]^x[227]^x[226]^x[188]^x[184]^x[183]^x[182]^x[173]^x[172]^x[171]^x[161]^x[119]^x[112]^x[109]^x[106]^x[98]^x[55]^x[43]^x[28]^x[24]^x[23]^x[18]^x[17]^x[13]^x[7];
	y[22]=x[346]^x[335]^x[283]^x[278]^x[272]^x[268]^x[257]^x[246]^x[237]^x[226]^x[225]^x[187]^x[183]^x[182]^x[181]^x[172]^x[171]^x[170]^x[160]^x[118]^x[111]^x[108]^x[105]^x[97]^x[54]^x[42]^x[27]^x[23]^x[22]^x[17]^x[16]^x[12]^x[6];
	y[21]=x[345]^x[334]^x[282]^x[277]^x[271]^x[267]^x[256]^x[245]^x[236]^x[225]^x[224]^x[186]^x[182]^x[181]^x[180]^x[171]^x[169]^x[117]^x[110]^x[107]^x[104]^x[96]^x[53]^x[41]^x[26]^x[22]^x[21]^x[16]^x[15]^x[11]^x[5];
	y[20]=x[287]^x[281]^x[276]^x[270]^x[255]^x[244]^x[235]^x[234]^x[224]^x[190]^x[181]^x[180]^x[170]^x[168]^x[127]^x[116]^x[52]^x[40]^x[21]^x[20]^x[15]^x[14]^x[10]^x[4];
	y[19]=x[286]^x[280]^x[275]^x[269]^x[255]^x[254]^x[243]^x[233]^x[189]^x[180]^x[179]^x[169]^x[167]^x[126]^x[115]^x[51]^x[39]^x[20]^x[19]^x[14]^x[13]^x[9]^x[3];
	y[18]=x[285]^x[279]^x[274]^x[268]^x[254]^x[253]^x[242]^x[232]^x[188]^x[179]^x[178]^x[168]^x[166]^x[125]^x[114]^x[50]^x[38]^x[19]^x[18]^x[13]^x[12]^x[8]^x[2];
	y[17]=x[341]^x[330]^x[284]^x[278]^x[273]^x[267]^x[253]^x[252]^x[241]^x[231]^x[187]^x[178]^x[177]^x[167]^x[165]^x[124]^x[113]^x[106]^x[100]^x[49]^x[37]^x[18]^x[17]^x[12]^x[11]^x[7]^x[1];
	y[16]=x[340]^x[329]^x[283]^x[277]^x[272]^x[266]^x[252]^x[251]^x[240]^x[230]^x[186]^x[177]^x[176]^x[166]^x[164]^x[123]^x[112]^x[105]^x[99]^x[48]^x[36]^x[17]^x[16]^x[11]^x[10]^x[6]^x[0];
	y[15]=x[339]^x[328]^x[282]^x[276]^x[271]^x[265]^x[251]^x[250]^x[239]^x[229]^x[185]^x[176]^x[175]^x[165]^x[163]^x[122]^x[111]^x[104]^x[98]^x[47]^x[35]^x[16]^x[15]^x[10]^x[9]^x[5];
	y[14]=x[338]^x[327]^x[281]^x[275]^x[270]^x[264]^x[250]^x[249]^x[238]^x[228]^x[184]^x[175]^x[174]^x[164]^x[162]^x[121]^x[110]^x[103]^x[97]^x[46]^x[34]^x[15]^x[14]^x[9]^x[8]^x[4];
	y[13]=x[337]^x[326]^x[280]^x[274]^x[269]^x[263]^x[249]^x[248]^x[237]^x[227]^x[183]^x[174]^x[173]^x[163]^x[161]^x[120]^x[109]^x[102]^x[96]^x[45]^x[33]^x[14]^x[13]^x[8]^x[7]^x[3];
	y[12]=x[336]^x[325]^x[279]^x[273]^x[268]^x[262]^x[248]^x[247]^x[236]^x[226]^x[182]^x[173]^x[172]^x[162]^x[160]^x[119]^x[108]^x[101]^x[44]^x[32]^x[13]^x[12]^x[7]^x[6]^x[2];
	y[11]=x[278]^x[272]^x[267]^x[261]^x[247]^x[246]^x[235]^x[225]^x[172]^x[171]^x[161]^x[118]^x[107]^x[43]^x[12]^x[11]^x[6]^x[5]^x[1];
	y[10]=x[277]^x[271]^x[266]^x[260]^x[246]^x[245]^x[234]^x[224]^x[171]^x[170]^x[160]^x[117]^x[106]^x[42]^x[11]^x[10]^x[5]^x[4]^x[0];
	y[9]=x[276]^x[270]^x[265]^x[259]^x[255]^x[245]^x[244]^x[234]^x[233]^x[191]^x[169]^x[116]^x[105]^x[41]^x[31]^x[25]^x[9]^x[3];
	y[8]=x[275]^x[269]^x[264]^x[258]^x[254]^x[244]^x[243]^x[233]^x[232]^x[190]^x[168]^x[115]^x[104]^x[40]^x[30]^x[24]^x[8]^x[2];
	y[7]=x[274]^x[268]^x[263]^x[257]^x[253]^x[243]^x[242]^x[232]^x[231]^x[189]^x[167]^x[114]^x[103]^x[39]^x[29]^x[23]^x[7]^x[1];
	y[6]=x[273]^x[267]^x[262]^x[256]^x[252]^x[242]^x[241]^x[231]^x[230]^x[188]^x[166]^x[113]^x[102]^x[38]^x[28]^x[22]^x[6]^x[0];
	y[5]=x[272]^x[261]^x[251]^x[241]^x[240]^x[230]^x[229]^x[187]^x[181]^x[175]^x[170]^x[165]^x[164]^x[112]^x[101]^x[37]^x[27]^x[10]^x[5];
	y[4]=x[271]^x[260]^x[250]^x[240]^x[239]^x[229]^x[228]^x[186]^x[180]^x[174]^x[169]^x[164]^x[163]^x[111]^x[100]^x[36]^x[26]^x[9]^x[4];
	y[3]=x[270]^x[259]^x[249]^x[239]^x[238]^x[228]^x[227]^x[185]^x[179]^x[173]^x[168]^x[163]^x[162]^x[110]^x[99]^x[35]^x[25]^x[8]^x[3];
	y[2]=x[269]^x[258]^x[248]^x[238]^x[237]^x[227]^x[226]^x[184]^x[178]^x[172]^x[167]^x[162]^x[161]^x[109]^x[98]^x[34]^x[24]^x[7]^x[2];
	y[1]=x[268]^x[257]^x[247]^x[237]^x[236]^x[226]^x[225]^x[183]^x[177]^x[171]^x[166]^x[161]^x[160]^x[108]^x[97]^x[33]^x[23]^x[6]^x[1];
	y[0]=x[267]^x[256]^x[246]^x[236]^x[235]^x[225]^x[224]^x[182]^x[176]^x[165]^x[160]^x[107]^x[96]^x[32]^x[22]^x[5]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint29(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[378]^x[377]^x[374]^x[368]^x[363]^x[362]^x[357]^x[356]^x[255]^x[249]^x[245]^x[242]^x[239]^x[236]^x[234]^x[231]^x[228]^x[225]^x[223]^x[214]^x[203]^x[202]^x[148]^x[95]^x[85]^x[82]^x[74]^x[71]^x[31]^x[19]^x[7];
	y[30]=x[382]^x[376]^x[373]^x[367]^x[362]^x[361]^x[356]^x[355]^x[254]^x[248]^x[244]^x[241]^x[238]^x[235]^x[233]^x[230]^x[227]^x[224]^x[222]^x[213]^x[202]^x[201]^x[94]^x[84]^x[81]^x[73]^x[70]^x[30]^x[18]^x[6];
	y[29]=x[381]^x[375]^x[372]^x[366]^x[361]^x[360]^x[355]^x[354]^x[253]^x[247]^x[243]^x[240]^x[237]^x[232]^x[229]^x[226]^x[221]^x[212]^x[201]^x[200]^x[93]^x[83]^x[80]^x[72]^x[69]^x[29]^x[17]^x[5];
	y[28]=x[380]^x[374]^x[371]^x[365]^x[360]^x[359]^x[354]^x[353]^x[252]^x[246]^x[242]^x[239]^x[236]^x[231]^x[228]^x[225]^x[220]^x[211]^x[200]^x[199]^x[92]^x[82]^x[79]^x[71]^x[68]^x[28]^x[16]^x[4];
	y[27]=x[379]^x[373]^x[370]^x[364]^x[359]^x[358]^x[353]^x[352]^x[251]^x[245]^x[241]^x[238]^x[235]^x[230]^x[227]^x[224]^x[219]^x[210]^x[199]^x[198]^x[91]^x[81]^x[78]^x[70]^x[67]^x[27]^x[15]^x[3];
	y[26]=x[378]^x[373]^x[372]^x[369]^x[363]^x[358]^x[357]^x[352]^x[318]^x[307]^x[255]^x[250]^x[244]^x[240]^x[237]^x[229]^x[226]^x[218]^x[209]^x[198]^x[197]^x[90]^x[83]^x[80]^x[69]^x[66]^x[26]^x[14]^x[2];
	y[25]=x[383]^x[377]^x[372]^x[371]^x[368]^x[357]^x[356]^x[317]^x[306]^x[254]^x[249]^x[243]^x[239]^x[236]^x[228]^x[225]^x[217]^x[208]^x[197]^x[196]^x[89]^x[82]^x[79]^x[68]^x[65]^x[25]^x[13]^x[1];
	y[24]=x[382]^x[376]^x[371]^x[370]^x[367]^x[356]^x[355]^x[316]^x[305]^x[253]^x[248]^x[242]^x[238]^x[235]^x[227]^x[224]^x[216]^x[207]^x[196]^x[195]^x[88]^x[81]^x[78]^x[67]^x[64]^x[24]^x[12]^x[0];
	y[23]=x[381]^x[375]^x[370]^x[369]^x[366]^x[355]^x[354]^x[315]^x[304]^x[252]^x[247]^x[241]^x[237]^x[226]^x[215]^x[206]^x[195]^x[194]^x[87]^x[80]^x[77]^x[74]^x[66]^x[23]^x[11];
	y[22]=x[380]^x[374]^x[369]^x[368]^x[365]^x[354]^x[353]^x[314]^x[303]^x[251]^x[246]^x[240]^x[236]^x[225]^x[214]^x[205]^x[194]^x[193]^x[86]^x[79]^x[76]^x[73]^x[65]^x[22]^x[10];
	y[21]=x[379]^x[373]^x[368]^x[367]^x[364]^x[353]^x[352]^x[313]^x[302]^x[250]^x[245]^x[239]^x[235]^x[224]^x[213]^x[204]^x[193]^x[192]^x[138]^x[85]^x[78]^x[75]^x[72]^x[64]^x[21]^x[9];
	y[20]=x[383]^x[378]^x[377]^x[372]^x[366]^x[363]^x[362]^x[356]^x[352]^x[255]^x[249]^x[244]^x[238]^x[223]^x[212]^x[203]^x[202]^x[192]^x[158]^x[137]^x[95]^x[84]^x[20]^x[8];
	y[19]=x[383]^x[382]^x[377]^x[376]^x[371]^x[365]^x[361]^x[355]^x[254]^x[248]^x[243]^x[237]^x[223]^x[222]^x[211]^x[201]^x[157]^x[136]^x[94]^x[83]^x[19]^x[7];
	y[18]=x[382]^x[381]^x[376]^x[375]^x[370]^x[364]^x[360]^x[354]^x[253]^x[247]^x[242]^x[236]^x[222]^x[221]^x[210]^x[200]^x[156]^x[135]^x[93]^x[82]^x[18]^x[6];
	y[17]=x[381]^x[380]^x[375]^x[374]^x[369]^x[363]^x[359]^x[353]^x[309]^x[298]^x[252]^x[246]^x[241]^x[235]^x[221]^x[220]^x[209]^x[199]^x[155]^x[134]^x[92]^x[81]^x[74]^x[68]^x[17]^x[5];
	y[16]=x[380]^x[379]^x[374]^x[373]^x[368]^x[362]^x[358]^x[352]^x[308]^x[297]^x[251]^x[245]^x[240]^x[234]^x[220]^x[219]^x[208]^x[198]^x[154]^x[133]^x[91]^x[80]^x[73]^x[67]^x[16]^x[4];
	y[15]=x[379]^x[378]^x[373]^x[372]^x[367]^x[362]^x[361]^x[357]^x[307]^x[296]^x[250]^x[244]^x[239]^x[233]^x[219]^x[218]^x[207]^x[197]^x[153]^x[132]^x[90]^x[79]^x[72]^x[66]^x[15]^x[3];
	y[14]=x[378]^x[377]^x[372]^x[371]^x[366]^x[361]^x[360]^x[356]^x[306]^x[295]^x[249]^x[243]^x[238]^x[232]^x[218]^x[217]^x[206]^x[196]^x[152]^x[131]^x[89]^x[78]^x[71]^x[65]^x[14]^x[2];
	y[13]=x[377]^x[376]^x[371]^x[370]^x[365]^x[360]^x[359]^x[355]^x[305]^x[294]^x[248]^x[242]^x[237]^x[231]^x[217]^x[216]^x[205]^x[195]^x[151]^x[130]^x[88]^x[77]^x[70]^x[64]^x[13]^x[1];
	y[12]=x[376]^x[375]^x[370]^x[369]^x[364]^x[359]^x[358]^x[354]^x[304]^x[293]^x[247]^x[241]^x[236]^x[230]^x[216]^x[215]^x[204]^x[194]^x[150]^x[129]^x[87]^x[76]^x[69]^x[12]^x[0];
	y[11]=x[375]^x[374]^x[369]^x[368]^x[363]^x[358]^x[357]^x[353]^x[246]^x[240]^x[235]^x[229]^x[215]^x[214]^x[203]^x[193]^x[128]^x[86]^x[75]^x[11];
	y[10]=x[374]^x[373]^x[368]^x[367]^x[362]^x[357]^x[356]^x[352]^x[245]^x[239]^x[234]^x[228]^x[214]^x[213]^x[202]^x[192]^x[85]^x[74]^x[10];
	y[9]=x[383]^x[377]^x[373]^x[372]^x[367]^x[366]^x[362]^x[361]^x[356]^x[355]^x[244]^x[238]^x[233]^x[227]^x[223]^x[213]^x[212]^x[202]^x[201]^x[147]^x[84]^x[73]^x[9];
	y[8]=x[382]^x[376]^x[372]^x[371]^x[366]^x[365]^x[361]^x[360]^x[355]^x[354]^x[243]^x[237]^x[232]^x[226]^x[222]^x[212]^x[211]^x[201]^x[200]^x[146]^x[83]^x[72]^x[8];
	y[7]=x[381]^x[375]^x[371]^x[370]^x[365]^x[364]^x[360]^x[359]^x[354]^x[353]^x[242]^x[236]^x[231]^x[225]^x[221]^x[211]^x[210]^x[200]^x[199]^x[145]^x[82]^x[71]^x[7];
	y[6]=x[380]^x[374]^x[370]^x[369]^x[364]^x[363]^x[359]^x[358]^x[353]^x[352]^x[241]^x[235]^x[230]^x[224]^x[220]^x[210]^x[209]^x[199]^x[198]^x[144]^x[81]^x[70]^x[6];
	y[5]=x[379]^x[373]^x[369]^x[368]^x[362]^x[358]^x[357]^x[240]^x[229]^x[219]^x[209]^x[208]^x[198]^x[197]^x[143]^x[80]^x[69]^x[5];
	y[4]=x[378]^x[372]^x[368]^x[367]^x[361]^x[357]^x[356]^x[239]^x[228]^x[218]^x[208]^x[207]^x[197]^x[196]^x[142]^x[79]^x[68]^x[4];
	y[3]=x[377]^x[371]^x[367]^x[366]^x[360]^x[356]^x[355]^x[238]^x[227]^x[217]^x[207]^x[206]^x[196]^x[195]^x[141]^x[78]^x[67]^x[3];
	y[2]=x[376]^x[370]^x[366]^x[365]^x[359]^x[355]^x[354]^x[237]^x[226]^x[216]^x[206]^x[205]^x[195]^x[194]^x[140]^x[77]^x[66]^x[2];
	y[1]=x[375]^x[369]^x[365]^x[364]^x[358]^x[354]^x[353]^x[236]^x[225]^x[215]^x[205]^x[204]^x[194]^x[193]^x[139]^x[76]^x[65]^x[1];
	y[0]=x[374]^x[368]^x[364]^x[363]^x[357]^x[353]^x[352]^x[235]^x[224]^x[214]^x[204]^x[203]^x[193]^x[192]^x[75]^x[64]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint30(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[373]^x[371]^x[370]^x[362]^x[359]^x[351]^x[346]^x[345]^x[342]^x[336]^x[331]^x[330]^x[325]^x[324]^x[223]^x[217]^x[213]^x[210]^x[207]^x[204]^x[202]^x[199]^x[196]^x[193]^x[191]^x[182]^x[171]^x[170]^x[159]^x[153]^x[147]^x[141]^x[135]^x[129]^x[116]^x[63]^x[53]^x[50]^x[42]^x[39];
	y[30]=x[382]^x[381]^x[372]^x[370]^x[369]^x[361]^x[358]^x[350]^x[344]^x[341]^x[335]^x[330]^x[329]^x[324]^x[323]^x[222]^x[216]^x[212]^x[209]^x[206]^x[203]^x[201]^x[198]^x[195]^x[192]^x[190]^x[181]^x[170]^x[169]^x[158]^x[152]^x[146]^x[140]^x[134]^x[128]^x[62]^x[52]^x[49]^x[41]^x[38];
	y[29]=x[381]^x[380]^x[371]^x[369]^x[368]^x[360]^x[357]^x[349]^x[343]^x[340]^x[334]^x[329]^x[328]^x[323]^x[322]^x[221]^x[215]^x[211]^x[208]^x[205]^x[200]^x[197]^x[194]^x[189]^x[180]^x[169]^x[168]^x[157]^x[151]^x[145]^x[139]^x[133]^x[61]^x[51]^x[48]^x[40]^x[37];
	y[28]=x[380]^x[379]^x[370]^x[368]^x[367]^x[359]^x[356]^x[348]^x[342]^x[339]^x[333]^x[328]^x[327]^x[322]^x[321]^x[220]^x[214]^x[210]^x[207]^x[204]^x[199]^x[196]^x[193]^x[188]^x[179]^x[168]^x[167]^x[156]^x[150]^x[144]^x[138]^x[132]^x[60]^x[50]^x[47]^x[39]^x[36];
	y[27]=x[379]^x[378]^x[369]^x[367]^x[366]^x[358]^x[355]^x[347]^x[341]^x[338]^x[332]^x[327]^x[326]^x[321]^x[320]^x[219]^x[213]^x[209]^x[206]^x[203]^x[198]^x[195]^x[192]^x[187]^x[178]^x[167]^x[166]^x[155]^x[149]^x[143]^x[137]^x[131]^x[59]^x[49]^x[46]^x[38]^x[35];
	y[26]=x[378]^x[377]^x[368]^x[366]^x[365]^x[357]^x[354]^x[346]^x[341]^x[340]^x[337]^x[331]^x[326]^x[325]^x[320]^x[286]^x[275]^x[223]^x[218]^x[212]^x[208]^x[205]^x[197]^x[194]^x[186]^x[177]^x[166]^x[165]^x[154]^x[148]^x[142]^x[136]^x[130]^x[58]^x[51]^x[48]^x[37]^x[34];
	y[25]=x[377]^x[376]^x[367]^x[365]^x[364]^x[356]^x[353]^x[351]^x[345]^x[340]^x[339]^x[336]^x[325]^x[324]^x[285]^x[274]^x[222]^x[217]^x[211]^x[207]^x[204]^x[196]^x[193]^x[185]^x[176]^x[165]^x[164]^x[153]^x[147]^x[141]^x[135]^x[129]^x[57]^x[50]^x[47]^x[36]^x[33];
	y[24]=x[376]^x[375]^x[366]^x[364]^x[363]^x[355]^x[352]^x[350]^x[344]^x[339]^x[338]^x[335]^x[324]^x[323]^x[284]^x[273]^x[221]^x[216]^x[210]^x[206]^x[203]^x[195]^x[192]^x[184]^x[175]^x[164]^x[163]^x[152]^x[146]^x[140]^x[134]^x[128]^x[56]^x[49]^x[46]^x[35]^x[32];
	y[23]=x[375]^x[374]^x[365]^x[363]^x[354]^x[349]^x[343]^x[338]^x[337]^x[334]^x[323]^x[322]^x[283]^x[272]^x[220]^x[215]^x[209]^x[205]^x[194]^x[183]^x[174]^x[163]^x[162]^x[151]^x[145]^x[139]^x[133]^x[55]^x[48]^x[45]^x[42]^x[34];
	y[22]=x[374]^x[373]^x[364]^x[362]^x[353]^x[348]^x[342]^x[337]^x[336]^x[333]^x[322]^x[321]^x[282]^x[271]^x[219]^x[214]^x[208]^x[204]^x[193]^x[182]^x[173]^x[162]^x[161]^x[150]^x[144]^x[138]^x[132]^x[54]^x[47]^x[44]^x[41]^x[33];
	y[21]=x[373]^x[372]^x[363]^x[361]^x[352]^x[347]^x[341]^x[336]^x[335]^x[332]^x[321]^x[320]^x[281]^x[270]^x[218]^x[213]^x[207]^x[203]^x[192]^x[181]^x[172]^x[161]^x[160]^x[149]^x[143]^x[137]^x[131]^x[106]^x[53]^x[46]^x[43]^x[40]^x[32];
	y[20]=x[383]^x[372]^x[371]^x[360]^x[351]^x[346]^x[345]^x[340]^x[334]^x[331]^x[330]^x[324]^x[320]^x[223]^x[217]^x[212]^x[206]^x[191]^x[180]^x[171]^x[170]^x[160]^x[148]^x[142]^x[136]^x[130]^x[126]^x[105]^x[63]^x[52];
	y[19]=x[382]^x[371]^x[370]^x[359]^x[351]^x[350]^x[345]^x[344]^x[339]^x[333]^x[329]^x[323]^x[222]^x[216]^x[211]^x[205]^x[191]^x[190]^x[179]^x[169]^x[147]^x[141]^x[135]^x[129]^x[125]^x[104]^x[62]^x[51];
	y[18]=x[381]^x[370]^x[369]^x[358]^x[350]^x[349]^x[344]^x[343]^x[338]^x[332]^x[328]^x[322]^x[221]^x[215]^x[210]^x[204]^x[190]^x[189]^x[178]^x[168]^x[146]^x[140]^x[134]^x[128]^x[124]^x[103]^x[61]^x[50];
	y[17]=x[380]^x[369]^x[368]^x[357]^x[349]^x[348]^x[343]^x[342]^x[337]^x[331]^x[327]^x[321]^x[277]^x[266]^x[220]^x[214]^x[209]^x[203]^x[189]^x[188]^x[177]^x[167]^x[145]^x[139]^x[133]^x[123]^x[102]^x[60]^x[49]^x[42]^x[36];
	y[16]=x[379]^x[368]^x[367]^x[356]^x[348]^x[347]^x[342]^x[341]^x[336]^x[330]^x[326]^x[320]^x[276]^x[265]^x[219]^x[213]^x[208]^x[202]^x[188]^x[187]^x[176]^x[166]^x[144]^x[138]^x[132]^x[122]^x[101]^x[59]^x[48]^x[41]^x[35];
	y[15]=x[378]^x[367]^x[366]^x[355]^x[347]^x[346]^x[341]^x[340]^x[335]^x[330]^x[329]^x[325]^x[275]^x[264]^x[218]^x[212]^x[207]^x[201]^x[187]^x[186]^x[175]^x[165]^x[143]^x[137]^x[131]^x[121]^x[100]^x[58]^x[47]^x[40]^x[34];
	y[14]=x[377]^x[366]^x[365]^x[354]^x[346]^x[345]^x[340]^x[339]^x[334]^x[329]^x[328]^x[324]^x[274]^x[263]^x[217]^x[211]^x[206]^x[200]^x[186]^x[185]^x[174]^x[164]^x[142]^x[136]^x[130]^x[120]^x[99]^x[57]^x[46]^x[39]^x[33];
	y[13]=x[376]^x[365]^x[364]^x[353]^x[345]^x[344]^x[339]^x[338]^x[333]^x[328]^x[327]^x[323]^x[273]^x[262]^x[216]^x[210]^x[205]^x[199]^x[185]^x[184]^x[173]^x[163]^x[141]^x[135]^x[129]^x[119]^x[98]^x[56]^x[45]^x[38]^x[32];
	y[12]=x[375]^x[364]^x[363]^x[352]^x[344]^x[343]^x[338]^x[337]^x[332]^x[327]^x[326]^x[322]^x[272]^x[261]^x[215]^x[209]^x[204]^x[198]^x[184]^x[183]^x[172]^x[162]^x[140]^x[134]^x[128]^x[118]^x[97]^x[55]^x[44]^x[37];
	y[11]=x[374]^x[363]^x[343]^x[342]^x[337]^x[336]^x[331]^x[326]^x[325]^x[321]^x[214]^x[208]^x[203]^x[197]^x[183]^x[182]^x[171]^x[161]^x[139]^x[133]^x[96]^x[54]^x[43];
	y[10]=x[373]^x[362]^x[342]^x[341]^x[336]^x[335]^x[330]^x[325]^x[324]^x[320]^x[213]^x[207]^x[202]^x[196]^x[182]^x[181]^x[170]^x[160]^x[138]^x[132]^x[53]^x[42];
	y[9]=x[372]^x[361]^x[351]^x[345]^x[341]^x[340]^x[335]^x[334]^x[330]^x[329]^x[324]^x[323]^x[212]^x[206]^x[201]^x[195]^x[191]^x[181]^x[180]^x[170]^x[169]^x[137]^x[131]^x[115]^x[52]^x[41];
	y[8]=x[371]^x[360]^x[350]^x[344]^x[340]^x[339]^x[334]^x[333]^x[329]^x[328]^x[323]^x[322]^x[211]^x[205]^x[200]^x[194]^x[190]^x[180]^x[179]^x[169]^x[168]^x[136]^x[130]^x[114]^x[51]^x[40];
	y[7]=x[370]^x[359]^x[349]^x[343]^x[339]^x[338]^x[333]^x[332]^x[328]^x[327]^x[322]^x[321]^x[210]^x[204]^x[199]^x[193]^x[189]^x[179]^x[178]^x[168]^x[167]^x[135]^x[129]^x[113]^x[50]^x[39];
	y[6]=x[369]^x[358]^x[348]^x[342]^x[338]^x[337]^x[332]^x[331]^x[327]^x[326]^x[321]^x[320]^x[209]^x[203]^x[198]^x[192]^x[188]^x[178]^x[177]^x[167]^x[166]^x[134]^x[128]^x[112]^x[49]^x[38];
	y[5]=x[368]^x[357]^x[347]^x[341]^x[337]^x[336]^x[330]^x[326]^x[325]^x[208]^x[197]^x[187]^x[177]^x[176]^x[166]^x[165]^x[133]^x[111]^x[48]^x[37];
	y[4]=x[367]^x[356]^x[346]^x[340]^x[336]^x[335]^x[329]^x[325]^x[324]^x[207]^x[196]^x[186]^x[176]^x[175]^x[165]^x[164]^x[132]^x[110]^x[47]^x[36];
	y[3]=x[366]^x[355]^x[345]^x[339]^x[335]^x[334]^x[328]^x[324]^x[323]^x[206]^x[195]^x[185]^x[175]^x[174]^x[164]^x[163]^x[131]^x[109]^x[46]^x[35];
	y[2]=x[365]^x[354]^x[344]^x[338]^x[334]^x[333]^x[327]^x[323]^x[322]^x[205]^x[194]^x[184]^x[174]^x[173]^x[163]^x[162]^x[130]^x[108]^x[45]^x[34];
	y[1]=x[364]^x[353]^x[343]^x[337]^x[333]^x[332]^x[326]^x[322]^x[321]^x[204]^x[193]^x[183]^x[173]^x[172]^x[162]^x[161]^x[129]^x[107]^x[44]^x[33];
	y[0]=x[363]^x[352]^x[342]^x[336]^x[332]^x[331]^x[325]^x[321]^x[320]^x[203]^x[192]^x[182]^x[172]^x[171]^x[161]^x[160]^x[128]^x[43]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint31(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[350]^x[341]^x[339]^x[338]^x[330]^x[327]^x[319]^x[314]^x[313]^x[310]^x[304]^x[299]^x[298]^x[293]^x[292]^x[191]^x[185]^x[181]^x[178]^x[175]^x[172]^x[170]^x[167]^x[164]^x[161]^x[159]^x[150]^x[139]^x[138]^x[127]^x[121]^x[115]^x[109]^x[103]^x[97]^x[84]^x[31]^x[21]^x[18]^x[10]^x[7];
	y[30]=x[350]^x[349]^x[340]^x[338]^x[337]^x[329]^x[326]^x[318]^x[312]^x[309]^x[303]^x[298]^x[297]^x[292]^x[291]^x[190]^x[184]^x[180]^x[177]^x[174]^x[171]^x[169]^x[166]^x[163]^x[160]^x[158]^x[149]^x[138]^x[137]^x[126]^x[120]^x[114]^x[108]^x[102]^x[96]^x[30]^x[20]^x[17]^x[9]^x[6];
	y[29]=x[349]^x[348]^x[339]^x[337]^x[336]^x[328]^x[325]^x[317]^x[311]^x[308]^x[302]^x[297]^x[296]^x[291]^x[290]^x[189]^x[183]^x[179]^x[176]^x[173]^x[168]^x[165]^x[162]^x[157]^x[148]^x[137]^x[136]^x[125]^x[119]^x[113]^x[107]^x[101]^x[29]^x[19]^x[16]^x[8]^x[5];
	y[28]=x[348]^x[347]^x[338]^x[336]^x[335]^x[327]^x[324]^x[316]^x[310]^x[307]^x[301]^x[296]^x[295]^x[290]^x[289]^x[188]^x[182]^x[178]^x[175]^x[172]^x[167]^x[164]^x[161]^x[156]^x[147]^x[136]^x[135]^x[124]^x[118]^x[112]^x[106]^x[100]^x[28]^x[18]^x[15]^x[7]^x[4];
	y[27]=x[347]^x[346]^x[337]^x[335]^x[334]^x[326]^x[323]^x[315]^x[309]^x[306]^x[300]^x[295]^x[294]^x[289]^x[288]^x[187]^x[181]^x[177]^x[174]^x[171]^x[166]^x[163]^x[160]^x[155]^x[146]^x[135]^x[134]^x[123]^x[117]^x[111]^x[105]^x[99]^x[27]^x[17]^x[14]^x[6]^x[3];
	y[26]=x[346]^x[345]^x[336]^x[334]^x[333]^x[325]^x[322]^x[314]^x[309]^x[308]^x[305]^x[299]^x[294]^x[293]^x[288]^x[254]^x[243]^x[191]^x[186]^x[180]^x[176]^x[173]^x[165]^x[162]^x[154]^x[145]^x[134]^x[133]^x[122]^x[116]^x[110]^x[104]^x[98]^x[26]^x[19]^x[16]^x[5]^x[2];
	y[25]=x[345]^x[344]^x[335]^x[333]^x[332]^x[324]^x[321]^x[319]^x[313]^x[308]^x[307]^x[304]^x[293]^x[292]^x[253]^x[242]^x[190]^x[185]^x[179]^x[175]^x[172]^x[164]^x[161]^x[153]^x[144]^x[133]^x[132]^x[121]^x[115]^x[109]^x[103]^x[97]^x[25]^x[18]^x[15]^x[4]^x[1];
	y[24]=x[344]^x[343]^x[334]^x[332]^x[331]^x[323]^x[320]^x[318]^x[312]^x[307]^x[306]^x[303]^x[292]^x[291]^x[252]^x[241]^x[189]^x[184]^x[178]^x[174]^x[171]^x[163]^x[160]^x[152]^x[143]^x[132]^x[131]^x[120]^x[114]^x[108]^x[102]^x[96]^x[24]^x[17]^x[14]^x[3]^x[0];
	y[23]=x[343]^x[342]^x[333]^x[331]^x[322]^x[317]^x[311]^x[306]^x[305]^x[302]^x[291]^x[290]^x[251]^x[240]^x[188]^x[183]^x[177]^x[173]^x[162]^x[151]^x[142]^x[131]^x[130]^x[119]^x[113]^x[107]^x[101]^x[23]^x[16]^x[13]^x[10]^x[2];
	y[22]=x[342]^x[341]^x[332]^x[330]^x[321]^x[316]^x[310]^x[305]^x[304]^x[301]^x[290]^x[289]^x[250]^x[239]^x[187]^x[182]^x[176]^x[172]^x[161]^x[150]^x[141]^x[130]^x[129]^x[118]^x[112]^x[106]^x[100]^x[22]^x[15]^x[12]^x[9]^x[1];
	y[21]=x[341]^x[340]^x[331]^x[329]^x[320]^x[315]^x[309]^x[304]^x[303]^x[300]^x[289]^x[288]^x[249]^x[238]^x[186]^x[181]^x[175]^x[171]^x[160]^x[149]^x[140]^x[129]^x[128]^x[117]^x[111]^x[105]^x[99]^x[74]^x[21]^x[14]^x[11]^x[8]^x[0];
	y[20]=x[351]^x[340]^x[339]^x[328]^x[319]^x[314]^x[313]^x[308]^x[302]^x[299]^x[298]^x[292]^x[288]^x[191]^x[185]^x[180]^x[174]^x[159]^x[148]^x[139]^x[138]^x[128]^x[116]^x[110]^x[104]^x[98]^x[94]^x[73]^x[31]^x[20];
	y[19]=x[350]^x[339]^x[338]^x[327]^x[319]^x[318]^x[313]^x[312]^x[307]^x[301]^x[297]^x[291]^x[190]^x[184]^x[179]^x[173]^x[159]^x[158]^x[147]^x[137]^x[115]^x[109]^x[103]^x[97]^x[93]^x[72]^x[30]^x[19];
	y[18]=x[349]^x[338]^x[337]^x[326]^x[318]^x[317]^x[312]^x[311]^x[306]^x[300]^x[296]^x[290]^x[189]^x[183]^x[178]^x[172]^x[158]^x[157]^x[146]^x[136]^x[114]^x[108]^x[102]^x[96]^x[92]^x[71]^x[29]^x[18];
	y[17]=x[348]^x[337]^x[336]^x[325]^x[317]^x[316]^x[311]^x[310]^x[305]^x[299]^x[295]^x[289]^x[245]^x[234]^x[188]^x[182]^x[177]^x[171]^x[157]^x[156]^x[145]^x[135]^x[113]^x[107]^x[101]^x[91]^x[70]^x[28]^x[17]^x[10]^x[4];
	y[16]=x[347]^x[336]^x[335]^x[324]^x[316]^x[315]^x[310]^x[309]^x[304]^x[298]^x[294]^x[288]^x[244]^x[233]^x[187]^x[181]^x[176]^x[170]^x[156]^x[155]^x[144]^x[134]^x[112]^x[106]^x[100]^x[90]^x[69]^x[27]^x[16]^x[9]^x[3];
	y[15]=x[346]^x[335]^x[334]^x[323]^x[315]^x[314]^x[309]^x[308]^x[303]^x[298]^x[297]^x[293]^x[243]^x[232]^x[186]^x[180]^x[175]^x[169]^x[155]^x[154]^x[143]^x[133]^x[111]^x[105]^x[99]^x[89]^x[68]^x[26]^x[15]^x[8]^x[2];
	y[14]=x[345]^x[334]^x[333]^x[322]^x[314]^x[313]^x[308]^x[307]^x[302]^x[297]^x[296]^x[292]^x[242]^x[231]^x[185]^x[179]^x[174]^x[168]^x[154]^x[153]^x[142]^x[132]^x[110]^x[104]^x[98]^x[88]^x[67]^x[25]^x[14]^x[7]^x[1];
	y[13]=x[344]^x[333]^x[332]^x[321]^x[313]^x[312]^x[307]^x[306]^x[301]^x[296]^x[295]^x[291]^x[241]^x[230]^x[184]^x[178]^x[173]^x[167]^x[153]^x[152]^x[141]^x[131]^x[109]^x[103]^x[97]^x[87]^x[66]^x[24]^x[13]^x[6]^x[0];
	y[12]=x[343]^x[332]^x[331]^x[320]^x[312]^x[311]^x[306]^x[305]^x[300]^x[295]^x[294]^x[290]^x[240]^x[229]^x[183]^x[177]^x[172]^x[166]^x[152]^x[151]^x[140]^x[130]^x[108]^x[102]^x[96]^x[86]^x[65]^x[23]^x[12]^x[5];
	y[11]=x[342]^x[331]^x[311]^x[310]^x[305]^x[304]^x[299]^x[294]^x[293]^x[289]^x[182]^x[176]^x[171]^x[165]^x[151]^x[150]^x[139]^x[129]^x[107]^x[101]^x[64]^x[22]^x[11];
	y[10]=x[341]^x[330]^x[310]^x[309]^x[304]^x[303]^x[298]^x[293]^x[292]^x[288]^x[181]^x[175]^x[170]^x[164]^x[150]^x[149]^x[138]^x[128]^x[106]^x[100]^x[21]^x[10];
	y[9]=x[340]^x[329]^x[319]^x[313]^x[309]^x[308]^x[303]^x[302]^x[298]^x[297]^x[292]^x[291]^x[180]^x[174]^x[169]^x[163]^x[159]^x[149]^x[148]^x[138]^x[137]^x[105]^x[99]^x[83]^x[20]^x[9];
	y[8]=x[339]^x[328]^x[318]^x[312]^x[308]^x[307]^x[302]^x[301]^x[297]^x[296]^x[291]^x[290]^x[179]^x[173]^x[168]^x[162]^x[158]^x[148]^x[147]^x[137]^x[136]^x[104]^x[98]^x[82]^x[19]^x[8];
	y[7]=x[338]^x[327]^x[317]^x[311]^x[307]^x[306]^x[301]^x[300]^x[296]^x[295]^x[290]^x[289]^x[178]^x[172]^x[167]^x[161]^x[157]^x[147]^x[146]^x[136]^x[135]^x[103]^x[97]^x[81]^x[18]^x[7];
	y[6]=x[337]^x[326]^x[316]^x[310]^x[306]^x[305]^x[300]^x[299]^x[295]^x[294]^x[289]^x[288]^x[177]^x[171]^x[166]^x[160]^x[156]^x[146]^x[145]^x[135]^x[134]^x[102]^x[96]^x[80]^x[17]^x[6];
	y[5]=x[336]^x[325]^x[315]^x[309]^x[305]^x[304]^x[298]^x[294]^x[293]^x[176]^x[165]^x[155]^x[145]^x[144]^x[134]^x[133]^x[101]^x[79]^x[16]^x[5];
	y[4]=x[335]^x[324]^x[314]^x[308]^x[304]^x[303]^x[297]^x[293]^x[292]^x[175]^x[164]^x[154]^x[144]^x[143]^x[133]^x[132]^x[100]^x[78]^x[15]^x[4];
	y[3]=x[334]^x[323]^x[313]^x[307]^x[303]^x[302]^x[296]^x[292]^x[291]^x[174]^x[163]^x[153]^x[143]^x[142]^x[132]^x[131]^x[99]^x[77]^x[14]^x[3];
	y[2]=x[333]^x[322]^x[312]^x[306]^x[302]^x[301]^x[295]^x[291]^x[290]^x[173]^x[162]^x[152]^x[142]^x[141]^x[131]^x[130]^x[98]^x[76]^x[13]^x[2];
	y[1]=x[332]^x[321]^x[311]^x[305]^x[301]^x[300]^x[294]^x[290]^x[289]^x[172]^x[161]^x[151]^x[141]^x[140]^x[130]^x[129]^x[97]^x[75]^x[12]^x[1];
	y[0]=x[331]^x[320]^x[310]^x[304]^x[300]^x[299]^x[293]^x[289]^x[288]^x[171]^x[160]^x[150]^x[140]^x[139]^x[129]^x[128]^x[96]^x[11]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint32(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[381]^x[373]^x[363]^x[359]^x[352]^x[319]^x[318]^x[309]^x[307]^x[306]^x[298]^x[295]^x[287]^x[282]^x[281]^x[278]^x[272]^x[267]^x[266]^x[261]^x[260]^x[127]^x[118]^x[107]^x[106]^x[95]^x[89]^x[83]^x[77]^x[71]^x[65]^x[52];
	y[30]=x[383]^x[382]^x[380]^x[372]^x[358]^x[318]^x[317]^x[308]^x[306]^x[305]^x[297]^x[294]^x[286]^x[280]^x[277]^x[271]^x[266]^x[265]^x[260]^x[259]^x[126]^x[117]^x[106]^x[105]^x[94]^x[88]^x[82]^x[76]^x[70]^x[64];
	y[29]=x[382]^x[381]^x[379]^x[371]^x[357]^x[317]^x[316]^x[307]^x[305]^x[304]^x[296]^x[293]^x[285]^x[279]^x[276]^x[270]^x[265]^x[264]^x[259]^x[258]^x[138]^x[125]^x[116]^x[105]^x[104]^x[93]^x[87]^x[81]^x[75]^x[69];
	y[28]=x[381]^x[380]^x[378]^x[370]^x[356]^x[316]^x[315]^x[306]^x[304]^x[303]^x[295]^x[292]^x[284]^x[278]^x[275]^x[269]^x[264]^x[263]^x[258]^x[257]^x[137]^x[124]^x[115]^x[104]^x[103]^x[92]^x[86]^x[80]^x[74]^x[68];
	y[27]=x[380]^x[379]^x[377]^x[369]^x[355]^x[315]^x[314]^x[305]^x[303]^x[302]^x[294]^x[291]^x[283]^x[277]^x[274]^x[268]^x[263]^x[262]^x[257]^x[256]^x[136]^x[123]^x[114]^x[103]^x[102]^x[91]^x[85]^x[79]^x[73]^x[67];
	y[26]=x[382]^x[379]^x[378]^x[371]^x[368]^x[365]^x[354]^x[314]^x[313]^x[304]^x[302]^x[301]^x[293]^x[290]^x[282]^x[277]^x[276]^x[273]^x[267]^x[262]^x[261]^x[256]^x[222]^x[211]^x[159]^x[147]^x[138]^x[122]^x[113]^x[102]^x[101]^x[90]^x[84]^x[78]^x[72]^x[66];
	y[25]=x[381]^x[378]^x[377]^x[370]^x[367]^x[364]^x[353]^x[313]^x[312]^x[303]^x[301]^x[300]^x[292]^x[289]^x[287]^x[281]^x[276]^x[275]^x[272]^x[261]^x[260]^x[221]^x[210]^x[158]^x[146]^x[137]^x[121]^x[112]^x[101]^x[100]^x[89]^x[83]^x[77]^x[71]^x[65];
	y[24]=x[380]^x[377]^x[376]^x[369]^x[366]^x[363]^x[352]^x[312]^x[311]^x[302]^x[300]^x[299]^x[291]^x[288]^x[286]^x[280]^x[275]^x[274]^x[271]^x[260]^x[259]^x[220]^x[209]^x[157]^x[145]^x[136]^x[120]^x[111]^x[100]^x[99]^x[88]^x[82]^x[76]^x[70]^x[64];
	y[23]=x[379]^x[376]^x[375]^x[373]^x[368]^x[365]^x[362]^x[311]^x[310]^x[301]^x[299]^x[290]^x[285]^x[279]^x[274]^x[273]^x[270]^x[259]^x[258]^x[219]^x[208]^x[156]^x[144]^x[135]^x[132]^x[119]^x[110]^x[99]^x[98]^x[87]^x[81]^x[75]^x[69];
	y[22]=x[378]^x[375]^x[374]^x[372]^x[367]^x[364]^x[361]^x[310]^x[309]^x[300]^x[298]^x[289]^x[284]^x[278]^x[273]^x[272]^x[269]^x[258]^x[257]^x[218]^x[207]^x[155]^x[143]^x[134]^x[131]^x[118]^x[109]^x[98]^x[97]^x[86]^x[80]^x[74]^x[68];
	y[21]=x[377]^x[374]^x[373]^x[371]^x[366]^x[363]^x[360]^x[309]^x[308]^x[299]^x[297]^x[288]^x[283]^x[277]^x[272]^x[271]^x[268]^x[257]^x[256]^x[217]^x[206]^x[154]^x[142]^x[133]^x[130]^x[117]^x[108]^x[97]^x[96]^x[85]^x[79]^x[73]^x[67]^x[42];
	y[20]=x[373]^x[372]^x[362]^x[319]^x[308]^x[307]^x[296]^x[287]^x[282]^x[281]^x[276]^x[270]^x[267]^x[266]^x[260]^x[256]^x[127]^x[116]^x[107]^x[106]^x[96]^x[84]^x[78]^x[72]^x[66]^x[62]^x[41];
	y[19]=x[372]^x[371]^x[361]^x[318]^x[307]^x[306]^x[295]^x[287]^x[286]^x[281]^x[280]^x[275]^x[269]^x[265]^x[259]^x[127]^x[126]^x[115]^x[105]^x[83]^x[77]^x[71]^x[65]^x[61]^x[40];
	y[18]=x[371]^x[370]^x[360]^x[317]^x[306]^x[305]^x[294]^x[286]^x[285]^x[280]^x[279]^x[274]^x[268]^x[264]^x[258]^x[126]^x[125]^x[114]^x[104]^x[82]^x[76]^x[70]^x[64]^x[60]^x[39];
	y[17]=x[373]^x[370]^x[369]^x[367]^x[362]^x[359]^x[356]^x[316]^x[305]^x[304]^x[293]^x[285]^x[284]^x[279]^x[278]^x[273]^x[267]^x[263]^x[257]^x[213]^x[202]^x[138]^x[125]^x[124]^x[113]^x[103]^x[81]^x[75]^x[69]^x[59]^x[38];
	y[16]=x[372]^x[369]^x[368]^x[366]^x[361]^x[358]^x[355]^x[315]^x[304]^x[303]^x[292]^x[284]^x[283]^x[278]^x[277]^x[272]^x[266]^x[262]^x[256]^x[212]^x[201]^x[137]^x[124]^x[123]^x[112]^x[102]^x[80]^x[74]^x[68]^x[58]^x[37];
	y[15]=x[371]^x[368]^x[367]^x[365]^x[360]^x[357]^x[354]^x[314]^x[303]^x[302]^x[291]^x[283]^x[282]^x[277]^x[276]^x[271]^x[266]^x[265]^x[261]^x[211]^x[200]^x[136]^x[123]^x[122]^x[111]^x[101]^x[79]^x[73]^x[67]^x[57]^x[36];
	y[14]=x[370]^x[367]^x[366]^x[364]^x[359]^x[356]^x[353]^x[313]^x[302]^x[301]^x[290]^x[282]^x[281]^x[276]^x[275]^x[270]^x[265]^x[264]^x[260]^x[210]^x[199]^x[135]^x[122]^x[121]^x[110]^x[100]^x[78]^x[72]^x[66]^x[56]^x[35];
	y[13]=x[369]^x[366]^x[365]^x[363]^x[358]^x[355]^x[352]^x[312]^x[301]^x[300]^x[289]^x[281]^x[280]^x[275]^x[274]^x[269]^x[264]^x[263]^x[259]^x[209]^x[198]^x[134]^x[121]^x[120]^x[109]^x[99]^x[77]^x[71]^x[65]^x[55]^x[34];
	y[12]=x[368]^x[365]^x[364]^x[357]^x[354]^x[311]^x[300]^x[299]^x[288]^x[280]^x[279]^x[274]^x[273]^x[268]^x[263]^x[262]^x[258]^x[208]^x[197]^x[133]^x[120]^x[119]^x[108]^x[98]^x[76]^x[70]^x[64]^x[54]^x[33];
	y[11]=x[364]^x[363]^x[353]^x[310]^x[299]^x[279]^x[278]^x[273]^x[272]^x[267]^x[262]^x[261]^x[257]^x[119]^x[118]^x[107]^x[97]^x[75]^x[69]^x[32];
	y[10]=x[363]^x[362]^x[352]^x[309]^x[298]^x[278]^x[277]^x[272]^x[271]^x[266]^x[261]^x[260]^x[256]^x[118]^x[117]^x[106]^x[96]^x[74]^x[68];
	y[9]=x[383]^x[361]^x[308]^x[297]^x[287]^x[281]^x[277]^x[276]^x[271]^x[270]^x[266]^x[265]^x[260]^x[259]^x[127]^x[117]^x[116]^x[106]^x[105]^x[73]^x[67]^x[51];
	y[8]=x[382]^x[360]^x[307]^x[296]^x[286]^x[280]^x[276]^x[275]^x[270]^x[269]^x[265]^x[264]^x[259]^x[258]^x[126]^x[116]^x[115]^x[105]^x[104]^x[72]^x[66]^x[50];
	y[7]=x[381]^x[359]^x[306]^x[295]^x[285]^x[279]^x[275]^x[274]^x[269]^x[268]^x[264]^x[263]^x[258]^x[257]^x[125]^x[115]^x[114]^x[104]^x[103]^x[71]^x[65]^x[49];
	y[6]=x[380]^x[358]^x[305]^x[294]^x[284]^x[278]^x[274]^x[273]^x[268]^x[267]^x[263]^x[262]^x[257]^x[256]^x[124]^x[114]^x[113]^x[103]^x[102]^x[70]^x[64]^x[48];
	y[5]=x[379]^x[357]^x[304]^x[293]^x[283]^x[277]^x[273]^x[272]^x[266]^x[262]^x[261]^x[138]^x[123]^x[113]^x[112]^x[102]^x[101]^x[69]^x[47];
	y[4]=x[378]^x[356]^x[303]^x[292]^x[282]^x[276]^x[272]^x[271]^x[265]^x[261]^x[260]^x[137]^x[122]^x[112]^x[111]^x[101]^x[100]^x[68]^x[46];
	y[3]=x[377]^x[355]^x[302]^x[291]^x[281]^x[275]^x[271]^x[270]^x[264]^x[260]^x[259]^x[136]^x[121]^x[111]^x[110]^x[100]^x[99]^x[67]^x[45];
	y[2]=x[376]^x[354]^x[301]^x[290]^x[280]^x[274]^x[270]^x[269]^x[263]^x[259]^x[258]^x[135]^x[120]^x[110]^x[109]^x[99]^x[98]^x[66]^x[44];
	y[1]=x[375]^x[353]^x[300]^x[289]^x[279]^x[273]^x[269]^x[268]^x[262]^x[258]^x[257]^x[134]^x[119]^x[109]^x[108]^x[98]^x[97]^x[65]^x[43];
	y[0]=x[374]^x[352]^x[299]^x[288]^x[278]^x[272]^x[268]^x[267]^x[261]^x[257]^x[256]^x[133]^x[118]^x[108]^x[107]^x[97]^x[96]^x[64];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint33(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[349]^x[341]^x[331]^x[327]^x[320]^x[287]^x[286]^x[277]^x[275]^x[274]^x[266]^x[263]^x[255]^x[250]^x[249]^x[246]^x[240]^x[235]^x[234]^x[229]^x[228]^x[95]^x[86]^x[75]^x[74]^x[63]^x[57]^x[51]^x[45]^x[39]^x[33]^x[20];
	y[30]=x[351]^x[350]^x[348]^x[340]^x[326]^x[286]^x[285]^x[276]^x[274]^x[273]^x[265]^x[262]^x[254]^x[248]^x[245]^x[239]^x[234]^x[233]^x[228]^x[227]^x[94]^x[85]^x[74]^x[73]^x[62]^x[56]^x[50]^x[44]^x[38]^x[32];
	y[29]=x[350]^x[349]^x[347]^x[339]^x[325]^x[285]^x[284]^x[275]^x[273]^x[272]^x[264]^x[261]^x[253]^x[247]^x[244]^x[238]^x[233]^x[232]^x[227]^x[226]^x[106]^x[93]^x[84]^x[73]^x[72]^x[61]^x[55]^x[49]^x[43]^x[37];
	y[28]=x[349]^x[348]^x[346]^x[338]^x[324]^x[284]^x[283]^x[274]^x[272]^x[271]^x[263]^x[260]^x[252]^x[246]^x[243]^x[237]^x[232]^x[231]^x[226]^x[225]^x[105]^x[92]^x[83]^x[72]^x[71]^x[60]^x[54]^x[48]^x[42]^x[36];
	y[27]=x[348]^x[347]^x[345]^x[337]^x[323]^x[283]^x[282]^x[273]^x[271]^x[270]^x[262]^x[259]^x[251]^x[245]^x[242]^x[236]^x[231]^x[230]^x[225]^x[224]^x[104]^x[91]^x[82]^x[71]^x[70]^x[59]^x[53]^x[47]^x[41]^x[35];
	y[26]=x[350]^x[347]^x[346]^x[339]^x[336]^x[333]^x[322]^x[282]^x[281]^x[272]^x[270]^x[269]^x[261]^x[258]^x[250]^x[245]^x[244]^x[241]^x[235]^x[230]^x[229]^x[224]^x[190]^x[179]^x[127]^x[115]^x[106]^x[90]^x[81]^x[70]^x[69]^x[58]^x[52]^x[46]^x[40]^x[34];
	y[25]=x[349]^x[346]^x[345]^x[338]^x[335]^x[332]^x[321]^x[281]^x[280]^x[271]^x[269]^x[268]^x[260]^x[257]^x[255]^x[249]^x[244]^x[243]^x[240]^x[229]^x[228]^x[189]^x[178]^x[126]^x[114]^x[105]^x[89]^x[80]^x[69]^x[68]^x[57]^x[51]^x[45]^x[39]^x[33];
	y[24]=x[348]^x[345]^x[344]^x[337]^x[334]^x[331]^x[320]^x[280]^x[279]^x[270]^x[268]^x[267]^x[259]^x[256]^x[254]^x[248]^x[243]^x[242]^x[239]^x[228]^x[227]^x[188]^x[177]^x[125]^x[113]^x[104]^x[88]^x[79]^x[68]^x[67]^x[56]^x[50]^x[44]^x[38]^x[32];
	y[23]=x[347]^x[344]^x[343]^x[341]^x[336]^x[333]^x[330]^x[279]^x[278]^x[269]^x[267]^x[258]^x[253]^x[247]^x[242]^x[241]^x[238]^x[227]^x[226]^x[187]^x[176]^x[124]^x[112]^x[103]^x[100]^x[87]^x[78]^x[67]^x[66]^x[55]^x[49]^x[43]^x[37];
	y[22]=x[346]^x[343]^x[342]^x[340]^x[335]^x[332]^x[329]^x[278]^x[277]^x[268]^x[266]^x[257]^x[252]^x[246]^x[241]^x[240]^x[237]^x[226]^x[225]^x[186]^x[175]^x[123]^x[111]^x[102]^x[99]^x[86]^x[77]^x[66]^x[65]^x[54]^x[48]^x[42]^x[36];
	y[21]=x[345]^x[342]^x[341]^x[339]^x[334]^x[331]^x[328]^x[277]^x[276]^x[267]^x[265]^x[256]^x[251]^x[245]^x[240]^x[239]^x[236]^x[225]^x[224]^x[185]^x[174]^x[122]^x[110]^x[101]^x[98]^x[85]^x[76]^x[65]^x[64]^x[53]^x[47]^x[41]^x[35]^x[10];
	y[20]=x[341]^x[340]^x[330]^x[287]^x[276]^x[275]^x[264]^x[255]^x[250]^x[249]^x[244]^x[238]^x[235]^x[234]^x[228]^x[224]^x[95]^x[84]^x[75]^x[74]^x[64]^x[52]^x[46]^x[40]^x[34]^x[30]^x[9];
	y[19]=x[340]^x[339]^x[329]^x[286]^x[275]^x[274]^x[263]^x[255]^x[254]^x[249]^x[248]^x[243]^x[237]^x[233]^x[227]^x[95]^x[94]^x[83]^x[73]^x[51]^x[45]^x[39]^x[33]^x[29]^x[8];
	y[18]=x[339]^x[338]^x[328]^x[285]^x[274]^x[273]^x[262]^x[254]^x[253]^x[248]^x[247]^x[242]^x[236]^x[232]^x[226]^x[94]^x[93]^x[82]^x[72]^x[50]^x[44]^x[38]^x[32]^x[28]^x[7];
	y[17]=x[341]^x[338]^x[337]^x[335]^x[330]^x[327]^x[324]^x[284]^x[273]^x[272]^x[261]^x[253]^x[252]^x[247]^x[246]^x[241]^x[235]^x[231]^x[225]^x[181]^x[170]^x[106]^x[93]^x[92]^x[81]^x[71]^x[49]^x[43]^x[37]^x[27]^x[6];
	y[16]=x[340]^x[337]^x[336]^x[334]^x[329]^x[326]^x[323]^x[283]^x[272]^x[271]^x[260]^x[252]^x[251]^x[246]^x[245]^x[240]^x[234]^x[230]^x[224]^x[180]^x[169]^x[105]^x[92]^x[91]^x[80]^x[70]^x[48]^x[42]^x[36]^x[26]^x[5];
	y[15]=x[339]^x[336]^x[335]^x[333]^x[328]^x[325]^x[322]^x[282]^x[271]^x[270]^x[259]^x[251]^x[250]^x[245]^x[244]^x[239]^x[234]^x[233]^x[229]^x[179]^x[168]^x[104]^x[91]^x[90]^x[79]^x[69]^x[47]^x[41]^x[35]^x[25]^x[4];
	y[14]=x[338]^x[335]^x[334]^x[332]^x[327]^x[324]^x[321]^x[281]^x[270]^x[269]^x[258]^x[250]^x[249]^x[244]^x[243]^x[238]^x[233]^x[232]^x[228]^x[178]^x[167]^x[103]^x[90]^x[89]^x[78]^x[68]^x[46]^x[40]^x[34]^x[24]^x[3];
	y[13]=x[337]^x[334]^x[333]^x[331]^x[326]^x[323]^x[320]^x[280]^x[269]^x[268]^x[257]^x[249]^x[248]^x[243]^x[242]^x[237]^x[232]^x[231]^x[227]^x[177]^x[166]^x[102]^x[89]^x[88]^x[77]^x[67]^x[45]^x[39]^x[33]^x[23]^x[2];
	y[12]=x[336]^x[333]^x[332]^x[325]^x[322]^x[279]^x[268]^x[267]^x[256]^x[248]^x[247]^x[242]^x[241]^x[236]^x[231]^x[230]^x[226]^x[176]^x[165]^x[101]^x[88]^x[87]^x[76]^x[66]^x[44]^x[38]^x[32]^x[22]^x[1];
	y[11]=x[332]^x[331]^x[321]^x[278]^x[267]^x[247]^x[246]^x[241]^x[240]^x[235]^x[230]^x[229]^x[225]^x[87]^x[86]^x[75]^x[65]^x[43]^x[37]^x[0];
	y[10]=x[331]^x[330]^x[320]^x[277]^x[266]^x[246]^x[245]^x[240]^x[239]^x[234]^x[229]^x[228]^x[224]^x[86]^x[85]^x[74]^x[64]^x[42]^x[36];
	y[9]=x[351]^x[329]^x[276]^x[265]^x[255]^x[249]^x[245]^x[244]^x[239]^x[238]^x[234]^x[233]^x[228]^x[227]^x[95]^x[85]^x[84]^x[74]^x[73]^x[41]^x[35]^x[19];
	y[8]=x[350]^x[328]^x[275]^x[264]^x[254]^x[248]^x[244]^x[243]^x[238]^x[237]^x[233]^x[232]^x[227]^x[226]^x[94]^x[84]^x[83]^x[73]^x[72]^x[40]^x[34]^x[18];
	y[7]=x[349]^x[327]^x[274]^x[263]^x[253]^x[247]^x[243]^x[242]^x[237]^x[236]^x[232]^x[231]^x[226]^x[225]^x[93]^x[83]^x[82]^x[72]^x[71]^x[39]^x[33]^x[17];
	y[6]=x[348]^x[326]^x[273]^x[262]^x[252]^x[246]^x[242]^x[241]^x[236]^x[235]^x[231]^x[230]^x[225]^x[224]^x[92]^x[82]^x[81]^x[71]^x[70]^x[38]^x[32]^x[16];
	y[5]=x[347]^x[325]^x[272]^x[261]^x[251]^x[245]^x[241]^x[240]^x[234]^x[230]^x[229]^x[106]^x[91]^x[81]^x[80]^x[70]^x[69]^x[37]^x[15];
	y[4]=x[346]^x[324]^x[271]^x[260]^x[250]^x[244]^x[240]^x[239]^x[233]^x[229]^x[228]^x[105]^x[90]^x[80]^x[79]^x[69]^x[68]^x[36]^x[14];
	y[3]=x[345]^x[323]^x[270]^x[259]^x[249]^x[243]^x[239]^x[238]^x[232]^x[228]^x[227]^x[104]^x[89]^x[79]^x[78]^x[68]^x[67]^x[35]^x[13];
	y[2]=x[344]^x[322]^x[269]^x[258]^x[248]^x[242]^x[238]^x[237]^x[231]^x[227]^x[226]^x[103]^x[88]^x[78]^x[77]^x[67]^x[66]^x[34]^x[12];
	y[1]=x[343]^x[321]^x[268]^x[257]^x[247]^x[241]^x[237]^x[236]^x[230]^x[226]^x[225]^x[102]^x[87]^x[77]^x[76]^x[66]^x[65]^x[33]^x[11];
	y[0]=x[342]^x[320]^x[267]^x[256]^x[246]^x[240]^x[236]^x[235]^x[229]^x[225]^x[224]^x[101]^x[86]^x[76]^x[75]^x[65]^x[64]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint34(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[372]^x[319]^x[317]^x[309]^x[299]^x[295]^x[288]^x[255]^x[254]^x[245]^x[243]^x[242]^x[234]^x[231]^x[223]^x[218]^x[217]^x[214]^x[208]^x[203]^x[202]^x[197]^x[196]^x[148]^x[142]^x[63]^x[54]^x[43]^x[42]^x[31]^x[25]^x[19]^x[13]^x[7]^x[1];
	y[30]=x[319]^x[318]^x[316]^x[308]^x[294]^x[254]^x[253]^x[244]^x[242]^x[241]^x[233]^x[230]^x[222]^x[216]^x[213]^x[207]^x[202]^x[201]^x[196]^x[195]^x[62]^x[53]^x[42]^x[41]^x[30]^x[24]^x[18]^x[12]^x[6]^x[0];
	y[29]=x[318]^x[317]^x[315]^x[307]^x[293]^x[253]^x[252]^x[243]^x[241]^x[240]^x[232]^x[229]^x[221]^x[215]^x[212]^x[206]^x[201]^x[200]^x[195]^x[194]^x[74]^x[61]^x[52]^x[41]^x[40]^x[29]^x[23]^x[17]^x[11]^x[5];
	y[28]=x[317]^x[316]^x[314]^x[306]^x[292]^x[252]^x[251]^x[242]^x[240]^x[239]^x[231]^x[228]^x[220]^x[214]^x[211]^x[205]^x[200]^x[199]^x[194]^x[193]^x[73]^x[60]^x[51]^x[40]^x[39]^x[28]^x[22]^x[16]^x[10]^x[4];
	y[27]=x[316]^x[315]^x[313]^x[305]^x[291]^x[251]^x[250]^x[241]^x[239]^x[238]^x[230]^x[227]^x[219]^x[213]^x[210]^x[204]^x[199]^x[198]^x[193]^x[192]^x[72]^x[59]^x[50]^x[39]^x[38]^x[27]^x[21]^x[15]^x[9]^x[3];
	y[26]=x[318]^x[315]^x[314]^x[307]^x[304]^x[301]^x[290]^x[250]^x[249]^x[240]^x[238]^x[237]^x[229]^x[226]^x[218]^x[213]^x[212]^x[209]^x[203]^x[198]^x[197]^x[192]^x[158]^x[147]^x[95]^x[83]^x[74]^x[58]^x[49]^x[38]^x[37]^x[26]^x[20]^x[14]^x[8]^x[2];
	y[25]=x[317]^x[314]^x[313]^x[306]^x[303]^x[300]^x[289]^x[249]^x[248]^x[239]^x[237]^x[236]^x[228]^x[225]^x[223]^x[217]^x[212]^x[211]^x[208]^x[197]^x[196]^x[157]^x[146]^x[94]^x[82]^x[73]^x[57]^x[48]^x[37]^x[36]^x[25]^x[19]^x[13]^x[7]^x[1];
	y[24]=x[316]^x[313]^x[312]^x[305]^x[302]^x[299]^x[288]^x[248]^x[247]^x[238]^x[236]^x[235]^x[227]^x[224]^x[222]^x[216]^x[211]^x[210]^x[207]^x[196]^x[195]^x[156]^x[145]^x[93]^x[81]^x[72]^x[56]^x[47]^x[36]^x[35]^x[24]^x[18]^x[12]^x[6]^x[0];
	y[23]=x[315]^x[312]^x[311]^x[309]^x[304]^x[301]^x[298]^x[247]^x[246]^x[237]^x[235]^x[226]^x[221]^x[215]^x[210]^x[209]^x[206]^x[195]^x[194]^x[155]^x[144]^x[92]^x[80]^x[71]^x[68]^x[55]^x[46]^x[35]^x[34]^x[23]^x[17]^x[11]^x[5];
	y[22]=x[314]^x[311]^x[310]^x[308]^x[303]^x[300]^x[297]^x[246]^x[245]^x[236]^x[234]^x[225]^x[220]^x[214]^x[209]^x[208]^x[205]^x[194]^x[193]^x[154]^x[143]^x[91]^x[79]^x[70]^x[67]^x[54]^x[45]^x[34]^x[33]^x[22]^x[16]^x[10]^x[4];
	y[21]=x[373]^x[362]^x[313]^x[310]^x[309]^x[307]^x[302]^x[299]^x[296]^x[245]^x[244]^x[235]^x[233]^x[224]^x[219]^x[213]^x[208]^x[207]^x[204]^x[193]^x[192]^x[153]^x[142]^x[138]^x[132]^x[90]^x[78]^x[69]^x[66]^x[53]^x[44]^x[33]^x[32]^x[21]^x[15]^x[9]^x[3];
	y[20]=x[382]^x[309]^x[308]^x[298]^x[255]^x[244]^x[243]^x[232]^x[223]^x[218]^x[217]^x[212]^x[206]^x[203]^x[202]^x[196]^x[192]^x[158]^x[152]^x[137]^x[131]^x[63]^x[52]^x[43]^x[42]^x[32]^x[20]^x[14]^x[8]^x[2];
	y[19]=x[381]^x[308]^x[307]^x[297]^x[254]^x[243]^x[242]^x[231]^x[223]^x[222]^x[217]^x[216]^x[211]^x[205]^x[201]^x[195]^x[157]^x[151]^x[136]^x[130]^x[63]^x[62]^x[51]^x[41]^x[19]^x[13]^x[7]^x[1];
	y[18]=x[380]^x[307]^x[306]^x[296]^x[253]^x[242]^x[241]^x[230]^x[222]^x[221]^x[216]^x[215]^x[210]^x[204]^x[200]^x[194]^x[156]^x[150]^x[135]^x[129]^x[62]^x[61]^x[50]^x[40]^x[18]^x[12]^x[6]^x[0];
	y[17]=x[379]^x[309]^x[306]^x[305]^x[303]^x[298]^x[295]^x[292]^x[252]^x[241]^x[240]^x[229]^x[221]^x[220]^x[215]^x[214]^x[209]^x[203]^x[199]^x[193]^x[155]^x[138]^x[134]^x[128]^x[74]^x[61]^x[60]^x[49]^x[39]^x[17]^x[11]^x[5];
	y[16]=x[378]^x[308]^x[305]^x[304]^x[302]^x[297]^x[294]^x[291]^x[251]^x[240]^x[239]^x[228]^x[220]^x[219]^x[214]^x[213]^x[208]^x[202]^x[198]^x[192]^x[154]^x[137]^x[133]^x[73]^x[60]^x[59]^x[48]^x[38]^x[16]^x[10]^x[4];
	y[15]=x[377]^x[307]^x[304]^x[303]^x[301]^x[296]^x[293]^x[290]^x[250]^x[239]^x[238]^x[227]^x[219]^x[218]^x[213]^x[212]^x[207]^x[202]^x[201]^x[197]^x[153]^x[136]^x[132]^x[72]^x[59]^x[58]^x[47]^x[37]^x[15]^x[9]^x[3];
	y[14]=x[376]^x[306]^x[303]^x[302]^x[300]^x[295]^x[292]^x[289]^x[249]^x[238]^x[237]^x[226]^x[218]^x[217]^x[212]^x[211]^x[206]^x[201]^x[200]^x[196]^x[152]^x[135]^x[131]^x[71]^x[58]^x[57]^x[46]^x[36]^x[14]^x[8]^x[2];
	y[13]=x[375]^x[305]^x[302]^x[301]^x[299]^x[294]^x[291]^x[288]^x[248]^x[237]^x[236]^x[225]^x[217]^x[216]^x[211]^x[210]^x[205]^x[200]^x[199]^x[195]^x[151]^x[134]^x[130]^x[70]^x[57]^x[56]^x[45]^x[35]^x[13]^x[7]^x[1];
	y[12]=x[374]^x[304]^x[301]^x[300]^x[293]^x[290]^x[247]^x[236]^x[235]^x[224]^x[216]^x[215]^x[210]^x[209]^x[204]^x[199]^x[198]^x[194]^x[150]^x[133]^x[129]^x[69]^x[56]^x[55]^x[44]^x[34]^x[12]^x[6]^x[0];
	y[11]=x[363]^x[352]^x[300]^x[299]^x[289]^x[246]^x[235]^x[215]^x[214]^x[209]^x[208]^x[203]^x[198]^x[197]^x[193]^x[128]^x[55]^x[54]^x[43]^x[33]^x[11]^x[5];
	y[10]=x[299]^x[298]^x[288]^x[245]^x[234]^x[214]^x[213]^x[208]^x[207]^x[202]^x[197]^x[196]^x[192]^x[54]^x[53]^x[42]^x[32]^x[10]^x[4];
	y[9]=x[382]^x[371]^x[319]^x[297]^x[244]^x[233]^x[223]^x[217]^x[213]^x[212]^x[207]^x[206]^x[202]^x[201]^x[196]^x[195]^x[147]^x[141]^x[63]^x[53]^x[52]^x[42]^x[41]^x[9]^x[3];
	y[8]=x[381]^x[370]^x[318]^x[296]^x[243]^x[232]^x[222]^x[216]^x[212]^x[211]^x[206]^x[205]^x[201]^x[200]^x[195]^x[194]^x[146]^x[140]^x[62]^x[52]^x[51]^x[41]^x[40]^x[8]^x[2];
	y[7]=x[380]^x[369]^x[317]^x[295]^x[242]^x[231]^x[221]^x[215]^x[211]^x[210]^x[205]^x[204]^x[200]^x[199]^x[194]^x[193]^x[145]^x[139]^x[61]^x[51]^x[50]^x[40]^x[39]^x[7]^x[1];
	y[6]=x[379]^x[368]^x[316]^x[294]^x[241]^x[230]^x[220]^x[214]^x[210]^x[209]^x[204]^x[203]^x[199]^x[198]^x[193]^x[192]^x[144]^x[138]^x[60]^x[50]^x[49]^x[39]^x[38]^x[6]^x[0];
	y[5]=x[378]^x[367]^x[315]^x[293]^x[240]^x[229]^x[219]^x[213]^x[209]^x[208]^x[202]^x[198]^x[197]^x[143]^x[137]^x[74]^x[59]^x[49]^x[48]^x[38]^x[37]^x[5];
	y[4]=x[377]^x[366]^x[314]^x[292]^x[239]^x[228]^x[218]^x[212]^x[208]^x[207]^x[201]^x[197]^x[196]^x[142]^x[136]^x[73]^x[58]^x[48]^x[47]^x[37]^x[36]^x[4];
	y[3]=x[376]^x[365]^x[313]^x[291]^x[238]^x[227]^x[217]^x[211]^x[207]^x[206]^x[200]^x[196]^x[195]^x[141]^x[135]^x[72]^x[57]^x[47]^x[46]^x[36]^x[35]^x[3];
	y[2]=x[375]^x[364]^x[312]^x[290]^x[237]^x[226]^x[216]^x[210]^x[206]^x[205]^x[199]^x[195]^x[194]^x[140]^x[134]^x[71]^x[56]^x[46]^x[45]^x[35]^x[34]^x[2];
	y[1]=x[374]^x[363]^x[311]^x[289]^x[236]^x[225]^x[215]^x[209]^x[205]^x[204]^x[198]^x[194]^x[193]^x[139]^x[133]^x[70]^x[55]^x[45]^x[44]^x[34]^x[33]^x[1];
	y[0]=x[310]^x[288]^x[235]^x[224]^x[214]^x[208]^x[204]^x[203]^x[197]^x[193]^x[192]^x[69]^x[54]^x[44]^x[43]^x[33]^x[32]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint35(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[377]^x[376]^x[373]^x[371]^x[370]^x[367]^x[365]^x[364]^x[362]^x[359]^x[356]^x[353]^x[351]^x[340]^x[287]^x[285]^x[277]^x[267]^x[263]^x[256]^x[223]^x[222]^x[213]^x[211]^x[210]^x[202]^x[199]^x[191]^x[186]^x[185]^x[182]^x[176]^x[171]^x[170]^x[165]^x[164]^x[159]^x[116]^x[110]^x[31]^x[22]^x[11]^x[10];
	y[30]=x[382]^x[381]^x[376]^x[375]^x[372]^x[370]^x[369]^x[366]^x[364]^x[363]^x[361]^x[358]^x[355]^x[352]^x[287]^x[286]^x[284]^x[276]^x[262]^x[222]^x[221]^x[212]^x[210]^x[209]^x[201]^x[198]^x[190]^x[184]^x[181]^x[175]^x[170]^x[169]^x[164]^x[163]^x[158]^x[30]^x[21]^x[10]^x[9];
	y[29]=x[381]^x[380]^x[375]^x[374]^x[371]^x[369]^x[368]^x[365]^x[363]^x[360]^x[357]^x[354]^x[286]^x[285]^x[283]^x[275]^x[261]^x[221]^x[220]^x[211]^x[209]^x[208]^x[200]^x[197]^x[189]^x[183]^x[180]^x[174]^x[169]^x[168]^x[163]^x[162]^x[157]^x[42]^x[29]^x[20]^x[9]^x[8];
	y[28]=x[380]^x[379]^x[374]^x[373]^x[370]^x[368]^x[367]^x[364]^x[362]^x[359]^x[356]^x[353]^x[285]^x[284]^x[282]^x[274]^x[260]^x[220]^x[219]^x[210]^x[208]^x[207]^x[199]^x[196]^x[188]^x[182]^x[179]^x[173]^x[168]^x[167]^x[162]^x[161]^x[156]^x[41]^x[28]^x[19]^x[8]^x[7];
	y[27]=x[379]^x[378]^x[373]^x[372]^x[369]^x[367]^x[366]^x[363]^x[361]^x[358]^x[355]^x[352]^x[284]^x[283]^x[281]^x[273]^x[259]^x[219]^x[218]^x[209]^x[207]^x[206]^x[198]^x[195]^x[187]^x[181]^x[178]^x[172]^x[167]^x[166]^x[161]^x[160]^x[155]^x[40]^x[27]^x[18]^x[7]^x[6];
	y[26]=x[383]^x[378]^x[377]^x[372]^x[371]^x[368]^x[366]^x[365]^x[360]^x[357]^x[354]^x[286]^x[283]^x[282]^x[275]^x[272]^x[269]^x[258]^x[218]^x[217]^x[208]^x[206]^x[205]^x[197]^x[194]^x[186]^x[181]^x[180]^x[177]^x[171]^x[166]^x[165]^x[160]^x[154]^x[126]^x[115]^x[63]^x[51]^x[42]^x[26]^x[17]^x[6]^x[5];
	y[25]=x[382]^x[377]^x[376]^x[371]^x[370]^x[367]^x[365]^x[364]^x[359]^x[356]^x[353]^x[285]^x[282]^x[281]^x[274]^x[271]^x[268]^x[257]^x[217]^x[216]^x[207]^x[205]^x[204]^x[196]^x[193]^x[191]^x[185]^x[180]^x[179]^x[176]^x[165]^x[164]^x[153]^x[125]^x[114]^x[62]^x[50]^x[41]^x[25]^x[16]^x[5]^x[4];
	y[24]=x[381]^x[376]^x[375]^x[370]^x[369]^x[366]^x[364]^x[363]^x[358]^x[355]^x[352]^x[284]^x[281]^x[280]^x[273]^x[270]^x[267]^x[256]^x[216]^x[215]^x[206]^x[204]^x[203]^x[195]^x[192]^x[190]^x[184]^x[179]^x[178]^x[175]^x[164]^x[163]^x[152]^x[124]^x[113]^x[61]^x[49]^x[40]^x[24]^x[15]^x[4]^x[3];
	y[23]=x[380]^x[375]^x[374]^x[369]^x[368]^x[365]^x[363]^x[357]^x[354]^x[283]^x[280]^x[279]^x[277]^x[272]^x[269]^x[266]^x[215]^x[214]^x[205]^x[203]^x[194]^x[189]^x[183]^x[178]^x[177]^x[174]^x[163]^x[162]^x[151]^x[123]^x[112]^x[60]^x[48]^x[39]^x[36]^x[23]^x[14]^x[3]^x[2];
	y[22]=x[379]^x[374]^x[373]^x[368]^x[367]^x[364]^x[362]^x[356]^x[353]^x[282]^x[279]^x[278]^x[276]^x[271]^x[268]^x[265]^x[214]^x[213]^x[204]^x[202]^x[193]^x[188]^x[182]^x[177]^x[176]^x[173]^x[162]^x[161]^x[150]^x[122]^x[111]^x[59]^x[47]^x[38]^x[35]^x[22]^x[13]^x[2]^x[1];
	y[21]=x[378]^x[373]^x[372]^x[367]^x[366]^x[363]^x[361]^x[355]^x[352]^x[341]^x[330]^x[281]^x[278]^x[277]^x[275]^x[270]^x[267]^x[264]^x[213]^x[212]^x[203]^x[201]^x[192]^x[187]^x[181]^x[176]^x[175]^x[172]^x[161]^x[160]^x[149]^x[121]^x[110]^x[106]^x[100]^x[58]^x[46]^x[37]^x[34]^x[21]^x[12]^x[1]^x[0];
	y[20]=x[383]^x[377]^x[372]^x[371]^x[366]^x[365]^x[360]^x[354]^x[350]^x[277]^x[276]^x[266]^x[223]^x[212]^x[211]^x[200]^x[191]^x[186]^x[185]^x[180]^x[174]^x[171]^x[170]^x[164]^x[160]^x[148]^x[126]^x[120]^x[105]^x[99]^x[31]^x[20]^x[11]^x[10]^x[0];
	y[19]=x[382]^x[376]^x[371]^x[370]^x[365]^x[364]^x[359]^x[353]^x[349]^x[276]^x[275]^x[265]^x[222]^x[211]^x[210]^x[199]^x[191]^x[190]^x[185]^x[184]^x[179]^x[173]^x[169]^x[163]^x[147]^x[125]^x[119]^x[104]^x[98]^x[31]^x[30]^x[19]^x[9];
	y[18]=x[381]^x[375]^x[370]^x[369]^x[364]^x[363]^x[358]^x[352]^x[348]^x[275]^x[274]^x[264]^x[221]^x[210]^x[209]^x[198]^x[190]^x[189]^x[184]^x[183]^x[178]^x[172]^x[168]^x[162]^x[146]^x[124]^x[118]^x[103]^x[97]^x[30]^x[29]^x[18]^x[8];
	y[17]=x[380]^x[374]^x[369]^x[368]^x[363]^x[357]^x[347]^x[277]^x[274]^x[273]^x[271]^x[266]^x[263]^x[260]^x[220]^x[209]^x[208]^x[197]^x[189]^x[188]^x[183]^x[182]^x[177]^x[171]^x[167]^x[161]^x[145]^x[123]^x[106]^x[102]^x[96]^x[42]^x[29]^x[28]^x[17]^x[7];
	y[16]=x[379]^x[373]^x[368]^x[367]^x[362]^x[356]^x[346]^x[276]^x[273]^x[272]^x[270]^x[265]^x[262]^x[259]^x[219]^x[208]^x[207]^x[196]^x[188]^x[187]^x[182]^x[181]^x[176]^x[170]^x[166]^x[160]^x[144]^x[122]^x[105]^x[101]^x[41]^x[28]^x[27]^x[16]^x[6];
	y[15]=x[378]^x[372]^x[367]^x[366]^x[361]^x[355]^x[345]^x[275]^x[272]^x[271]^x[269]^x[264]^x[261]^x[258]^x[218]^x[207]^x[206]^x[195]^x[187]^x[186]^x[181]^x[180]^x[175]^x[170]^x[169]^x[165]^x[143]^x[121]^x[104]^x[100]^x[40]^x[27]^x[26]^x[15]^x[5];
	y[14]=x[377]^x[371]^x[366]^x[365]^x[360]^x[354]^x[344]^x[274]^x[271]^x[270]^x[268]^x[263]^x[260]^x[257]^x[217]^x[206]^x[205]^x[194]^x[186]^x[185]^x[180]^x[179]^x[174]^x[169]^x[168]^x[164]^x[142]^x[120]^x[103]^x[99]^x[39]^x[26]^x[25]^x[14]^x[4];
	y[13]=x[376]^x[370]^x[365]^x[364]^x[359]^x[353]^x[343]^x[273]^x[270]^x[269]^x[267]^x[262]^x[259]^x[256]^x[216]^x[205]^x[204]^x[193]^x[185]^x[184]^x[179]^x[178]^x[173]^x[168]^x[167]^x[163]^x[141]^x[119]^x[102]^x[98]^x[38]^x[25]^x[24]^x[13]^x[3];
	y[12]=x[375]^x[369]^x[364]^x[363]^x[358]^x[352]^x[342]^x[272]^x[269]^x[268]^x[261]^x[258]^x[215]^x[204]^x[203]^x[192]^x[184]^x[183]^x[178]^x[177]^x[172]^x[167]^x[166]^x[162]^x[140]^x[118]^x[101]^x[97]^x[37]^x[24]^x[23]^x[12]^x[2];
	y[11]=x[374]^x[368]^x[363]^x[357]^x[331]^x[320]^x[268]^x[267]^x[257]^x[214]^x[203]^x[183]^x[182]^x[177]^x[176]^x[171]^x[166]^x[165]^x[161]^x[139]^x[96]^x[23]^x[22]^x[11]^x[1];
	y[10]=x[373]^x[367]^x[362]^x[356]^x[267]^x[266]^x[256]^x[213]^x[202]^x[182]^x[181]^x[176]^x[175]^x[170]^x[165]^x[164]^x[160]^x[138]^x[22]^x[21]^x[10]^x[0];
	y[9]=x[372]^x[366]^x[361]^x[355]^x[350]^x[339]^x[287]^x[265]^x[212]^x[201]^x[191]^x[185]^x[181]^x[180]^x[175]^x[174]^x[170]^x[169]^x[164]^x[163]^x[137]^x[115]^x[109]^x[31]^x[21]^x[20]^x[10]^x[9];
	y[8]=x[371]^x[365]^x[360]^x[354]^x[349]^x[338]^x[286]^x[264]^x[211]^x[200]^x[190]^x[184]^x[180]^x[179]^x[174]^x[173]^x[169]^x[168]^x[163]^x[162]^x[136]^x[114]^x[108]^x[30]^x[20]^x[19]^x[9]^x[8];
	y[7]=x[370]^x[364]^x[359]^x[353]^x[348]^x[337]^x[285]^x[263]^x[210]^x[199]^x[189]^x[183]^x[179]^x[178]^x[173]^x[172]^x[168]^x[167]^x[162]^x[161]^x[135]^x[113]^x[107]^x[29]^x[19]^x[18]^x[8]^x[7];
	y[6]=x[369]^x[363]^x[358]^x[352]^x[347]^x[336]^x[284]^x[262]^x[209]^x[198]^x[188]^x[182]^x[178]^x[177]^x[172]^x[171]^x[167]^x[166]^x[161]^x[160]^x[134]^x[112]^x[106]^x[28]^x[18]^x[17]^x[7]^x[6];
	y[5]=x[368]^x[357]^x[346]^x[335]^x[283]^x[261]^x[208]^x[197]^x[187]^x[181]^x[177]^x[176]^x[170]^x[166]^x[165]^x[133]^x[111]^x[105]^x[42]^x[27]^x[17]^x[16]^x[6]^x[5];
	y[4]=x[367]^x[356]^x[345]^x[334]^x[282]^x[260]^x[207]^x[196]^x[186]^x[180]^x[176]^x[175]^x[169]^x[165]^x[164]^x[132]^x[110]^x[104]^x[41]^x[26]^x[16]^x[15]^x[5]^x[4];
	y[3]=x[366]^x[355]^x[344]^x[333]^x[281]^x[259]^x[206]^x[195]^x[185]^x[179]^x[175]^x[174]^x[168]^x[164]^x[163]^x[131]^x[109]^x[103]^x[40]^x[25]^x[15]^x[14]^x[4]^x[3];
	y[2]=x[365]^x[354]^x[343]^x[332]^x[280]^x[258]^x[205]^x[194]^x[184]^x[178]^x[174]^x[173]^x[167]^x[163]^x[162]^x[130]^x[108]^x[102]^x[39]^x[24]^x[14]^x[13]^x[3]^x[2];
	y[1]=x[364]^x[353]^x[342]^x[331]^x[279]^x[257]^x[204]^x[193]^x[183]^x[177]^x[173]^x[172]^x[166]^x[162]^x[161]^x[129]^x[107]^x[101]^x[38]^x[23]^x[13]^x[12]^x[2]^x[1];
	y[0]=x[363]^x[352]^x[278]^x[256]^x[203]^x[192]^x[182]^x[176]^x[172]^x[171]^x[165]^x[161]^x[160]^x[128]^x[37]^x[22]^x[12]^x[11]^x[1]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint36(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[364]^x[363]^x[353]^x[351]^x[350]^x[345]^x[344]^x[341]^x[339]^x[338]^x[335]^x[333]^x[332]^x[330]^x[327]^x[324]^x[321]^x[319]^x[308]^x[255]^x[253]^x[245]^x[235]^x[231]^x[224]^x[191]^x[190]^x[181]^x[179]^x[178]^x[170]^x[167]^x[154]^x[127]^x[84]^x[78];
	y[30]=x[382]^x[363]^x[362]^x[352]^x[350]^x[349]^x[344]^x[343]^x[340]^x[338]^x[337]^x[334]^x[332]^x[331]^x[329]^x[326]^x[323]^x[320]^x[255]^x[254]^x[252]^x[244]^x[230]^x[190]^x[189]^x[180]^x[178]^x[177]^x[169]^x[166]^x[126];
	y[29]=x[383]^x[381]^x[361]^x[349]^x[348]^x[343]^x[342]^x[339]^x[337]^x[336]^x[333]^x[331]^x[328]^x[325]^x[322]^x[254]^x[253]^x[251]^x[243]^x[229]^x[189]^x[188]^x[179]^x[177]^x[176]^x[168]^x[165]^x[125]^x[10];
	y[28]=x[382]^x[380]^x[360]^x[348]^x[347]^x[342]^x[341]^x[338]^x[336]^x[335]^x[332]^x[330]^x[327]^x[324]^x[321]^x[253]^x[252]^x[250]^x[242]^x[228]^x[188]^x[187]^x[178]^x[176]^x[175]^x[167]^x[164]^x[124]^x[9];
	y[27]=x[381]^x[379]^x[359]^x[347]^x[346]^x[341]^x[340]^x[337]^x[335]^x[334]^x[331]^x[329]^x[326]^x[323]^x[320]^x[252]^x[251]^x[249]^x[241]^x[227]^x[187]^x[186]^x[177]^x[175]^x[174]^x[166]^x[163]^x[123]^x[8];
	y[26]=x[380]^x[378]^x[358]^x[351]^x[346]^x[345]^x[340]^x[339]^x[336]^x[334]^x[333]^x[328]^x[325]^x[322]^x[254]^x[251]^x[250]^x[243]^x[240]^x[237]^x[226]^x[186]^x[185]^x[176]^x[174]^x[173]^x[165]^x[162]^x[149]^x[122]^x[94]^x[83]^x[31]^x[19]^x[10];
	y[25]=x[379]^x[377]^x[357]^x[350]^x[345]^x[344]^x[339]^x[338]^x[335]^x[333]^x[332]^x[327]^x[324]^x[321]^x[253]^x[250]^x[249]^x[242]^x[239]^x[236]^x[225]^x[185]^x[184]^x[175]^x[173]^x[172]^x[164]^x[161]^x[159]^x[148]^x[138]^x[121]^x[93]^x[82]^x[30]^x[18]^x[9];
	y[24]=x[378]^x[376]^x[356]^x[349]^x[344]^x[343]^x[338]^x[337]^x[334]^x[332]^x[331]^x[326]^x[323]^x[320]^x[252]^x[249]^x[248]^x[241]^x[238]^x[235]^x[224]^x[184]^x[183]^x[174]^x[172]^x[171]^x[163]^x[160]^x[158]^x[147]^x[137]^x[120]^x[92]^x[81]^x[29]^x[17]^x[8];
	y[23]=x[377]^x[375]^x[355]^x[348]^x[343]^x[342]^x[337]^x[336]^x[333]^x[331]^x[325]^x[322]^x[251]^x[248]^x[247]^x[245]^x[240]^x[237]^x[234]^x[183]^x[182]^x[173]^x[171]^x[162]^x[157]^x[146]^x[136]^x[119]^x[91]^x[80]^x[28]^x[16]^x[7]^x[4];
	y[22]=x[376]^x[374]^x[354]^x[347]^x[342]^x[341]^x[336]^x[335]^x[332]^x[330]^x[324]^x[321]^x[250]^x[247]^x[246]^x[244]^x[239]^x[236]^x[233]^x[182]^x[181]^x[172]^x[170]^x[161]^x[156]^x[145]^x[135]^x[118]^x[90]^x[79]^x[27]^x[15]^x[6]^x[3];
	y[21]=x[375]^x[373]^x[353]^x[346]^x[341]^x[340]^x[335]^x[334]^x[331]^x[329]^x[323]^x[320]^x[309]^x[298]^x[249]^x[246]^x[245]^x[243]^x[238]^x[235]^x[232]^x[181]^x[180]^x[171]^x[169]^x[160]^x[155]^x[144]^x[134]^x[117]^x[89]^x[78]^x[74]^x[68]^x[26]^x[14]^x[5]^x[2];
	y[20]=x[374]^x[372]^x[352]^x[351]^x[345]^x[340]^x[339]^x[334]^x[333]^x[328]^x[322]^x[318]^x[245]^x[244]^x[234]^x[191]^x[180]^x[179]^x[168]^x[154]^x[133]^x[116]^x[94]^x[88]^x[73]^x[67];
	y[19]=x[383]^x[373]^x[371]^x[362]^x[350]^x[344]^x[339]^x[338]^x[333]^x[332]^x[327]^x[321]^x[317]^x[244]^x[243]^x[233]^x[190]^x[179]^x[178]^x[167]^x[115]^x[93]^x[87]^x[72]^x[66];
	y[18]=x[382]^x[372]^x[370]^x[361]^x[349]^x[343]^x[338]^x[337]^x[332]^x[331]^x[326]^x[320]^x[316]^x[243]^x[242]^x[232]^x[189]^x[178]^x[177]^x[166]^x[114]^x[92]^x[86]^x[71]^x[65];
	y[17]=x[381]^x[371]^x[369]^x[360]^x[348]^x[342]^x[337]^x[336]^x[331]^x[325]^x[315]^x[245]^x[242]^x[241]^x[239]^x[234]^x[231]^x[228]^x[188]^x[177]^x[176]^x[165]^x[113]^x[91]^x[74]^x[70]^x[64]^x[10];
	y[16]=x[380]^x[370]^x[368]^x[359]^x[347]^x[341]^x[336]^x[335]^x[330]^x[324]^x[314]^x[244]^x[241]^x[240]^x[238]^x[233]^x[230]^x[227]^x[187]^x[176]^x[175]^x[164]^x[112]^x[90]^x[73]^x[69]^x[9];
	y[15]=x[379]^x[369]^x[367]^x[358]^x[346]^x[340]^x[335]^x[334]^x[329]^x[323]^x[313]^x[243]^x[240]^x[239]^x[237]^x[232]^x[229]^x[226]^x[186]^x[175]^x[174]^x[163]^x[138]^x[111]^x[89]^x[72]^x[68]^x[8];
	y[14]=x[378]^x[368]^x[366]^x[357]^x[345]^x[339]^x[334]^x[333]^x[328]^x[322]^x[312]^x[242]^x[239]^x[238]^x[236]^x[231]^x[228]^x[225]^x[185]^x[174]^x[173]^x[162]^x[137]^x[110]^x[88]^x[71]^x[67]^x[7];
	y[13]=x[377]^x[367]^x[365]^x[356]^x[344]^x[338]^x[333]^x[332]^x[327]^x[321]^x[311]^x[241]^x[238]^x[237]^x[235]^x[230]^x[227]^x[224]^x[184]^x[173]^x[172]^x[161]^x[136]^x[109]^x[87]^x[70]^x[66]^x[6];
	y[12]=x[376]^x[366]^x[364]^x[355]^x[343]^x[337]^x[332]^x[331]^x[326]^x[320]^x[310]^x[240]^x[237]^x[236]^x[229]^x[226]^x[183]^x[172]^x[171]^x[160]^x[135]^x[108]^x[86]^x[69]^x[65]^x[5];
	y[11]=x[375]^x[365]^x[363]^x[354]^x[342]^x[336]^x[331]^x[325]^x[299]^x[288]^x[236]^x[235]^x[225]^x[182]^x[171]^x[134]^x[107]^x[64];
	y[10]=x[374]^x[364]^x[362]^x[353]^x[341]^x[335]^x[330]^x[324]^x[235]^x[234]^x[224]^x[181]^x[170]^x[133]^x[106];
	y[9]=x[373]^x[363]^x[361]^x[352]^x[340]^x[334]^x[329]^x[323]^x[318]^x[307]^x[255]^x[233]^x[180]^x[169]^x[105]^x[83]^x[77];
	y[8]=x[383]^x[372]^x[360]^x[339]^x[333]^x[328]^x[322]^x[317]^x[306]^x[254]^x[232]^x[179]^x[168]^x[104]^x[82]^x[76];
	y[7]=x[382]^x[371]^x[359]^x[338]^x[332]^x[327]^x[321]^x[316]^x[305]^x[253]^x[231]^x[178]^x[167]^x[103]^x[81]^x[75];
	y[6]=x[381]^x[370]^x[358]^x[337]^x[331]^x[326]^x[320]^x[315]^x[304]^x[252]^x[230]^x[177]^x[166]^x[102]^x[80]^x[74];
	y[5]=x[380]^x[369]^x[357]^x[336]^x[325]^x[314]^x[303]^x[251]^x[229]^x[176]^x[165]^x[139]^x[128]^x[101]^x[79]^x[73]^x[10];
	y[4]=x[379]^x[368]^x[356]^x[335]^x[324]^x[313]^x[302]^x[250]^x[228]^x[175]^x[164]^x[138]^x[100]^x[78]^x[72]^x[9];
	y[3]=x[378]^x[367]^x[355]^x[334]^x[323]^x[312]^x[301]^x[249]^x[227]^x[174]^x[163]^x[137]^x[99]^x[77]^x[71]^x[8];
	y[2]=x[377]^x[366]^x[354]^x[333]^x[322]^x[311]^x[300]^x[248]^x[226]^x[173]^x[162]^x[136]^x[98]^x[76]^x[70]^x[7];
	y[1]=x[376]^x[365]^x[353]^x[332]^x[321]^x[310]^x[299]^x[247]^x[225]^x[172]^x[161]^x[135]^x[97]^x[75]^x[69]^x[6];
	y[0]=x[375]^x[364]^x[352]^x[331]^x[320]^x[246]^x[224]^x[171]^x[160]^x[134]^x[96]^x[5];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint37(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[332]^x[331]^x[321]^x[319]^x[318]^x[313]^x[312]^x[309]^x[307]^x[306]^x[303]^x[301]^x[300]^x[298]^x[295]^x[292]^x[289]^x[287]^x[276]^x[223]^x[221]^x[213]^x[203]^x[199]^x[192]^x[159]^x[158]^x[149]^x[147]^x[146]^x[138]^x[135]^x[122]^x[95]^x[52]^x[46];
	y[30]=x[350]^x[331]^x[330]^x[320]^x[318]^x[317]^x[312]^x[311]^x[308]^x[306]^x[305]^x[302]^x[300]^x[299]^x[297]^x[294]^x[291]^x[288]^x[223]^x[222]^x[220]^x[212]^x[198]^x[158]^x[157]^x[148]^x[146]^x[145]^x[137]^x[134]^x[94];
	y[29]=x[373]^x[362]^x[351]^x[349]^x[329]^x[317]^x[316]^x[311]^x[310]^x[307]^x[305]^x[304]^x[301]^x[299]^x[296]^x[293]^x[290]^x[222]^x[221]^x[219]^x[211]^x[197]^x[157]^x[156]^x[147]^x[145]^x[144]^x[138]^x[136]^x[133]^x[132]^x[93];
	y[28]=x[372]^x[361]^x[350]^x[348]^x[328]^x[316]^x[315]^x[310]^x[309]^x[306]^x[304]^x[303]^x[300]^x[298]^x[295]^x[292]^x[289]^x[221]^x[220]^x[218]^x[210]^x[196]^x[156]^x[155]^x[146]^x[144]^x[143]^x[137]^x[135]^x[132]^x[131]^x[92];
	y[27]=x[371]^x[360]^x[349]^x[347]^x[327]^x[315]^x[314]^x[309]^x[308]^x[305]^x[303]^x[302]^x[299]^x[297]^x[294]^x[291]^x[288]^x[220]^x[219]^x[217]^x[209]^x[195]^x[155]^x[154]^x[145]^x[143]^x[142]^x[136]^x[134]^x[131]^x[130]^x[91];
	y[26]=x[383]^x[382]^x[371]^x[348]^x[346]^x[326]^x[319]^x[314]^x[313]^x[308]^x[307]^x[304]^x[302]^x[301]^x[296]^x[293]^x[290]^x[222]^x[219]^x[218]^x[211]^x[208]^x[205]^x[194]^x[159]^x[154]^x[147]^x[144]^x[142]^x[138]^x[133]^x[132]^x[130]^x[117]^x[90]^x[62]^x[51];
	y[25]=x[382]^x[381]^x[370]^x[347]^x[345]^x[325]^x[318]^x[313]^x[312]^x[307]^x[306]^x[303]^x[301]^x[300]^x[295]^x[292]^x[289]^x[221]^x[218]^x[217]^x[210]^x[207]^x[204]^x[193]^x[158]^x[153]^x[146]^x[143]^x[141]^x[137]^x[132]^x[131]^x[129]^x[127]^x[116]^x[106]^x[89]^x[61]^x[50];
	y[24]=x[381]^x[380]^x[369]^x[346]^x[344]^x[324]^x[317]^x[312]^x[311]^x[306]^x[305]^x[302]^x[300]^x[299]^x[294]^x[291]^x[288]^x[220]^x[217]^x[216]^x[209]^x[206]^x[203]^x[192]^x[157]^x[152]^x[145]^x[142]^x[140]^x[136]^x[131]^x[130]^x[128]^x[126]^x[115]^x[105]^x[88]^x[60]^x[49];
	y[23]=x[380]^x[379]^x[368]^x[367]^x[356]^x[345]^x[343]^x[323]^x[316]^x[311]^x[310]^x[305]^x[304]^x[301]^x[299]^x[293]^x[290]^x[219]^x[216]^x[215]^x[213]^x[208]^x[205]^x[202]^x[156]^x[151]^x[144]^x[141]^x[139]^x[138]^x[135]^x[132]^x[130]^x[129]^x[125]^x[114]^x[104]^x[87]^x[59]^x[48];
	y[22]=x[379]^x[378]^x[367]^x[366]^x[355]^x[344]^x[342]^x[322]^x[315]^x[310]^x[309]^x[304]^x[303]^x[300]^x[298]^x[292]^x[289]^x[218]^x[215]^x[214]^x[212]^x[207]^x[204]^x[201]^x[155]^x[150]^x[143]^x[140]^x[138]^x[137]^x[134]^x[131]^x[129]^x[128]^x[124]^x[113]^x[103]^x[86]^x[58]^x[47];
	y[21]=x[378]^x[377]^x[366]^x[365]^x[354]^x[343]^x[341]^x[321]^x[314]^x[309]^x[308]^x[303]^x[302]^x[299]^x[297]^x[291]^x[288]^x[277]^x[266]^x[217]^x[214]^x[213]^x[211]^x[206]^x[203]^x[200]^x[154]^x[149]^x[142]^x[139]^x[137]^x[136]^x[133]^x[130]^x[128]^x[123]^x[112]^x[102]^x[85]^x[57]^x[46]^x[42]^x[36];
	y[20]=x[342]^x[340]^x[320]^x[319]^x[313]^x[308]^x[307]^x[302]^x[301]^x[296]^x[290]^x[286]^x[213]^x[212]^x[202]^x[159]^x[148]^x[147]^x[136]^x[122]^x[101]^x[84]^x[62]^x[56]^x[41]^x[35];
	y[19]=x[351]^x[341]^x[339]^x[330]^x[318]^x[312]^x[307]^x[306]^x[301]^x[300]^x[295]^x[289]^x[285]^x[212]^x[211]^x[201]^x[158]^x[147]^x[146]^x[135]^x[83]^x[61]^x[55]^x[40]^x[34];
	y[18]=x[350]^x[340]^x[338]^x[329]^x[317]^x[311]^x[306]^x[305]^x[300]^x[299]^x[294]^x[288]^x[284]^x[211]^x[210]^x[200]^x[157]^x[146]^x[145]^x[134]^x[82]^x[60]^x[54]^x[39]^x[33];
	y[17]=x[373]^x[362]^x[349]^x[339]^x[337]^x[328]^x[316]^x[310]^x[305]^x[304]^x[299]^x[293]^x[283]^x[213]^x[210]^x[209]^x[207]^x[202]^x[199]^x[196]^x[156]^x[145]^x[144]^x[138]^x[133]^x[132]^x[81]^x[59]^x[42]^x[38]^x[32];
	y[16]=x[372]^x[361]^x[348]^x[338]^x[336]^x[327]^x[315]^x[309]^x[304]^x[303]^x[298]^x[292]^x[282]^x[212]^x[209]^x[208]^x[206]^x[201]^x[198]^x[195]^x[155]^x[144]^x[143]^x[137]^x[132]^x[131]^x[80]^x[58]^x[41]^x[37];
	y[15]=x[371]^x[360]^x[347]^x[337]^x[335]^x[326]^x[314]^x[308]^x[303]^x[302]^x[297]^x[291]^x[281]^x[211]^x[208]^x[207]^x[205]^x[200]^x[197]^x[194]^x[154]^x[143]^x[142]^x[136]^x[131]^x[130]^x[106]^x[79]^x[57]^x[40]^x[36];
	y[14]=x[370]^x[359]^x[346]^x[336]^x[334]^x[325]^x[313]^x[307]^x[302]^x[301]^x[296]^x[290]^x[280]^x[210]^x[207]^x[206]^x[204]^x[199]^x[196]^x[193]^x[153]^x[142]^x[141]^x[135]^x[130]^x[129]^x[105]^x[78]^x[56]^x[39]^x[35];
	y[13]=x[369]^x[358]^x[345]^x[335]^x[333]^x[324]^x[312]^x[306]^x[301]^x[300]^x[295]^x[289]^x[279]^x[209]^x[206]^x[205]^x[203]^x[198]^x[195]^x[192]^x[152]^x[141]^x[140]^x[134]^x[129]^x[128]^x[104]^x[77]^x[55]^x[38]^x[34];
	y[12]=x[368]^x[357]^x[344]^x[334]^x[332]^x[323]^x[311]^x[305]^x[300]^x[299]^x[294]^x[288]^x[278]^x[208]^x[205]^x[204]^x[197]^x[194]^x[151]^x[140]^x[139]^x[133]^x[128]^x[103]^x[76]^x[54]^x[37]^x[33];
	y[11]=x[343]^x[333]^x[331]^x[322]^x[310]^x[304]^x[299]^x[293]^x[267]^x[256]^x[204]^x[203]^x[193]^x[150]^x[139]^x[102]^x[75]^x[32];
	y[10]=x[342]^x[332]^x[330]^x[321]^x[309]^x[303]^x[298]^x[292]^x[203]^x[202]^x[192]^x[149]^x[138]^x[101]^x[74];
	y[9]=x[341]^x[331]^x[329]^x[320]^x[308]^x[302]^x[297]^x[291]^x[286]^x[275]^x[223]^x[201]^x[148]^x[137]^x[73]^x[51]^x[45];
	y[8]=x[351]^x[340]^x[328]^x[307]^x[301]^x[296]^x[290]^x[285]^x[274]^x[222]^x[200]^x[147]^x[136]^x[72]^x[50]^x[44];
	y[7]=x[350]^x[339]^x[327]^x[306]^x[300]^x[295]^x[289]^x[284]^x[273]^x[221]^x[199]^x[146]^x[135]^x[71]^x[49]^x[43];
	y[6]=x[349]^x[338]^x[326]^x[305]^x[299]^x[294]^x[288]^x[283]^x[272]^x[220]^x[198]^x[145]^x[134]^x[70]^x[48]^x[42];
	y[5]=x[373]^x[362]^x[348]^x[337]^x[325]^x[304]^x[293]^x[282]^x[271]^x[219]^x[197]^x[144]^x[138]^x[133]^x[132]^x[107]^x[96]^x[69]^x[47]^x[41];
	y[4]=x[372]^x[361]^x[347]^x[336]^x[324]^x[303]^x[292]^x[281]^x[270]^x[218]^x[196]^x[143]^x[137]^x[132]^x[131]^x[106]^x[68]^x[46]^x[40];
	y[3]=x[371]^x[360]^x[346]^x[335]^x[323]^x[302]^x[291]^x[280]^x[269]^x[217]^x[195]^x[142]^x[136]^x[131]^x[130]^x[105]^x[67]^x[45]^x[39];
	y[2]=x[370]^x[359]^x[345]^x[334]^x[322]^x[301]^x[290]^x[279]^x[268]^x[216]^x[194]^x[141]^x[135]^x[130]^x[129]^x[104]^x[66]^x[44]^x[38];
	y[1]=x[369]^x[358]^x[344]^x[333]^x[321]^x[300]^x[289]^x[278]^x[267]^x[215]^x[193]^x[140]^x[134]^x[129]^x[128]^x[103]^x[65]^x[43]^x[37];
	y[0]=x[368]^x[357]^x[343]^x[332]^x[320]^x[299]^x[288]^x[214]^x[192]^x[139]^x[133]^x[128]^x[102]^x[64];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint38(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[319]^x[300]^x[299]^x[289]^x[287]^x[286]^x[281]^x[280]^x[277]^x[275]^x[274]^x[271]^x[269]^x[268]^x[266]^x[263]^x[260]^x[257]^x[255]^x[244]^x[191]^x[189]^x[181]^x[171]^x[167]^x[160]^x[127]^x[126]^x[117]^x[115]^x[114]^x[106]^x[103]^x[90]^x[63]^x[20]^x[14];
	y[30]=x[318]^x[299]^x[298]^x[288]^x[286]^x[285]^x[280]^x[279]^x[276]^x[274]^x[273]^x[270]^x[268]^x[267]^x[265]^x[262]^x[259]^x[256]^x[191]^x[190]^x[188]^x[180]^x[166]^x[126]^x[125]^x[116]^x[114]^x[113]^x[105]^x[102]^x[62];
	y[29]=x[341]^x[330]^x[319]^x[317]^x[297]^x[285]^x[284]^x[279]^x[278]^x[275]^x[273]^x[272]^x[269]^x[267]^x[264]^x[261]^x[258]^x[190]^x[189]^x[187]^x[179]^x[165]^x[125]^x[124]^x[115]^x[113]^x[112]^x[106]^x[104]^x[101]^x[100]^x[61];
	y[28]=x[340]^x[329]^x[318]^x[316]^x[296]^x[284]^x[283]^x[278]^x[277]^x[274]^x[272]^x[271]^x[268]^x[266]^x[263]^x[260]^x[257]^x[189]^x[188]^x[186]^x[178]^x[164]^x[124]^x[123]^x[114]^x[112]^x[111]^x[105]^x[103]^x[100]^x[99]^x[60];
	y[27]=x[339]^x[328]^x[317]^x[315]^x[295]^x[283]^x[282]^x[277]^x[276]^x[273]^x[271]^x[270]^x[267]^x[265]^x[262]^x[259]^x[256]^x[188]^x[187]^x[185]^x[177]^x[163]^x[123]^x[122]^x[113]^x[111]^x[110]^x[104]^x[102]^x[99]^x[98]^x[59];
	y[26]=x[351]^x[350]^x[339]^x[316]^x[314]^x[294]^x[287]^x[282]^x[281]^x[276]^x[275]^x[272]^x[270]^x[269]^x[264]^x[261]^x[258]^x[190]^x[187]^x[186]^x[179]^x[176]^x[173]^x[162]^x[127]^x[122]^x[115]^x[112]^x[110]^x[106]^x[101]^x[100]^x[98]^x[85]^x[58]^x[30]^x[19];
	y[25]=x[350]^x[349]^x[338]^x[315]^x[313]^x[293]^x[286]^x[281]^x[280]^x[275]^x[274]^x[271]^x[269]^x[268]^x[263]^x[260]^x[257]^x[189]^x[186]^x[185]^x[178]^x[175]^x[172]^x[161]^x[126]^x[121]^x[114]^x[111]^x[109]^x[105]^x[100]^x[99]^x[97]^x[95]^x[84]^x[74]^x[57]^x[29]^x[18];
	y[24]=x[349]^x[348]^x[337]^x[314]^x[312]^x[292]^x[285]^x[280]^x[279]^x[274]^x[273]^x[270]^x[268]^x[267]^x[262]^x[259]^x[256]^x[188]^x[185]^x[184]^x[177]^x[174]^x[171]^x[160]^x[125]^x[120]^x[113]^x[110]^x[108]^x[104]^x[99]^x[98]^x[96]^x[94]^x[83]^x[73]^x[56]^x[28]^x[17];
	y[23]=x[348]^x[347]^x[336]^x[335]^x[324]^x[313]^x[311]^x[291]^x[284]^x[279]^x[278]^x[273]^x[272]^x[269]^x[267]^x[261]^x[258]^x[187]^x[184]^x[183]^x[181]^x[176]^x[173]^x[170]^x[124]^x[119]^x[112]^x[109]^x[107]^x[106]^x[103]^x[100]^x[98]^x[97]^x[93]^x[82]^x[72]^x[55]^x[27]^x[16];
	y[22]=x[347]^x[346]^x[335]^x[334]^x[323]^x[312]^x[310]^x[290]^x[283]^x[278]^x[277]^x[272]^x[271]^x[268]^x[266]^x[260]^x[257]^x[186]^x[183]^x[182]^x[180]^x[175]^x[172]^x[169]^x[123]^x[118]^x[111]^x[108]^x[106]^x[105]^x[102]^x[99]^x[97]^x[96]^x[92]^x[81]^x[71]^x[54]^x[26]^x[15];
	y[21]=x[346]^x[345]^x[334]^x[333]^x[322]^x[311]^x[309]^x[289]^x[282]^x[277]^x[276]^x[271]^x[270]^x[267]^x[265]^x[259]^x[256]^x[245]^x[234]^x[185]^x[182]^x[181]^x[179]^x[174]^x[171]^x[168]^x[122]^x[117]^x[110]^x[107]^x[105]^x[104]^x[101]^x[98]^x[96]^x[91]^x[80]^x[70]^x[53]^x[25]^x[14]^x[10]^x[4];
	y[20]=x[310]^x[308]^x[288]^x[287]^x[281]^x[276]^x[275]^x[270]^x[269]^x[264]^x[258]^x[254]^x[181]^x[180]^x[170]^x[127]^x[116]^x[115]^x[104]^x[90]^x[69]^x[52]^x[30]^x[24]^x[9]^x[3];
	y[19]=x[319]^x[309]^x[307]^x[298]^x[286]^x[280]^x[275]^x[274]^x[269]^x[268]^x[263]^x[257]^x[253]^x[180]^x[179]^x[169]^x[126]^x[115]^x[114]^x[103]^x[51]^x[29]^x[23]^x[8]^x[2];
	y[18]=x[318]^x[308]^x[306]^x[297]^x[285]^x[279]^x[274]^x[273]^x[268]^x[267]^x[262]^x[256]^x[252]^x[179]^x[178]^x[168]^x[125]^x[114]^x[113]^x[102]^x[50]^x[28]^x[22]^x[7]^x[1];
	y[17]=x[341]^x[330]^x[317]^x[307]^x[305]^x[296]^x[284]^x[278]^x[273]^x[272]^x[267]^x[261]^x[251]^x[181]^x[178]^x[177]^x[175]^x[170]^x[167]^x[164]^x[124]^x[113]^x[112]^x[106]^x[101]^x[100]^x[49]^x[27]^x[10]^x[6]^x[0];
	y[16]=x[340]^x[329]^x[316]^x[306]^x[304]^x[295]^x[283]^x[277]^x[272]^x[271]^x[266]^x[260]^x[250]^x[180]^x[177]^x[176]^x[174]^x[169]^x[166]^x[163]^x[123]^x[112]^x[111]^x[105]^x[100]^x[99]^x[48]^x[26]^x[9]^x[5];
	y[15]=x[339]^x[328]^x[315]^x[305]^x[303]^x[294]^x[282]^x[276]^x[271]^x[270]^x[265]^x[259]^x[249]^x[179]^x[176]^x[175]^x[173]^x[168]^x[165]^x[162]^x[122]^x[111]^x[110]^x[104]^x[99]^x[98]^x[74]^x[47]^x[25]^x[8]^x[4];
	y[14]=x[338]^x[327]^x[314]^x[304]^x[302]^x[293]^x[281]^x[275]^x[270]^x[269]^x[264]^x[258]^x[248]^x[178]^x[175]^x[174]^x[172]^x[167]^x[164]^x[161]^x[121]^x[110]^x[109]^x[103]^x[98]^x[97]^x[73]^x[46]^x[24]^x[7]^x[3];
	y[13]=x[337]^x[326]^x[313]^x[303]^x[301]^x[292]^x[280]^x[274]^x[269]^x[268]^x[263]^x[257]^x[247]^x[177]^x[174]^x[173]^x[171]^x[166]^x[163]^x[160]^x[120]^x[109]^x[108]^x[102]^x[97]^x[96]^x[72]^x[45]^x[23]^x[6]^x[2];
	y[12]=x[336]^x[325]^x[312]^x[302]^x[300]^x[291]^x[279]^x[273]^x[268]^x[267]^x[262]^x[256]^x[246]^x[176]^x[173]^x[172]^x[165]^x[162]^x[119]^x[108]^x[107]^x[101]^x[96]^x[71]^x[44]^x[22]^x[5]^x[1];
	y[11]=x[311]^x[301]^x[299]^x[290]^x[278]^x[272]^x[267]^x[261]^x[235]^x[224]^x[172]^x[171]^x[161]^x[118]^x[107]^x[70]^x[43]^x[0];
	y[10]=x[310]^x[300]^x[298]^x[289]^x[277]^x[271]^x[266]^x[260]^x[171]^x[170]^x[160]^x[117]^x[106]^x[69]^x[42];
	y[9]=x[309]^x[299]^x[297]^x[288]^x[276]^x[270]^x[265]^x[259]^x[254]^x[243]^x[191]^x[169]^x[116]^x[105]^x[41]^x[19]^x[13];
	y[8]=x[319]^x[308]^x[296]^x[275]^x[269]^x[264]^x[258]^x[253]^x[242]^x[190]^x[168]^x[115]^x[104]^x[40]^x[18]^x[12];
	y[7]=x[318]^x[307]^x[295]^x[274]^x[268]^x[263]^x[257]^x[252]^x[241]^x[189]^x[167]^x[114]^x[103]^x[39]^x[17]^x[11];
	y[6]=x[317]^x[306]^x[294]^x[273]^x[267]^x[262]^x[256]^x[251]^x[240]^x[188]^x[166]^x[113]^x[102]^x[38]^x[16]^x[10];
	y[5]=x[341]^x[330]^x[316]^x[305]^x[293]^x[272]^x[261]^x[250]^x[239]^x[187]^x[165]^x[112]^x[106]^x[101]^x[100]^x[75]^x[64]^x[37]^x[15]^x[9];
	y[4]=x[340]^x[329]^x[315]^x[304]^x[292]^x[271]^x[260]^x[249]^x[238]^x[186]^x[164]^x[111]^x[105]^x[100]^x[99]^x[74]^x[36]^x[14]^x[8];
	y[3]=x[339]^x[328]^x[314]^x[303]^x[291]^x[270]^x[259]^x[248]^x[237]^x[185]^x[163]^x[110]^x[104]^x[99]^x[98]^x[73]^x[35]^x[13]^x[7];
	y[2]=x[338]^x[327]^x[313]^x[302]^x[290]^x[269]^x[258]^x[247]^x[236]^x[184]^x[162]^x[109]^x[103]^x[98]^x[97]^x[72]^x[34]^x[12]^x[6];
	y[1]=x[337]^x[326]^x[312]^x[301]^x[289]^x[268]^x[257]^x[246]^x[235]^x[183]^x[161]^x[108]^x[102]^x[97]^x[96]^x[71]^x[33]^x[11]^x[5];
	y[0]=x[336]^x[325]^x[311]^x[300]^x[288]^x[267]^x[256]^x[182]^x[160]^x[107]^x[101]^x[96]^x[70]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint39(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[377]^x[372]^x[366]^x[287]^x[268]^x[267]^x[257]^x[255]^x[254]^x[249]^x[248]^x[245]^x[243]^x[242]^x[239]^x[237]^x[236]^x[234]^x[231]^x[228]^x[225]^x[223]^x[212]^x[159]^x[157]^x[149]^x[148]^x[139]^x[136]^x[135]^x[128]^x[95]^x[94]^x[85]^x[83]^x[82]^x[74]^x[71]^x[58]^x[31];
	y[30]=x[286]^x[267]^x[266]^x[256]^x[254]^x[253]^x[248]^x[247]^x[244]^x[242]^x[241]^x[238]^x[236]^x[235]^x[233]^x[230]^x[227]^x[224]^x[159]^x[158]^x[156]^x[148]^x[134]^x[94]^x[93]^x[84]^x[82]^x[81]^x[73]^x[70]^x[30];
	y[29]=x[309]^x[298]^x[287]^x[285]^x[265]^x[253]^x[252]^x[247]^x[246]^x[243]^x[241]^x[240]^x[237]^x[235]^x[232]^x[229]^x[226]^x[158]^x[157]^x[155]^x[147]^x[133]^x[93]^x[92]^x[83]^x[81]^x[80]^x[74]^x[72]^x[69]^x[68]^x[29];
	y[28]=x[308]^x[297]^x[286]^x[284]^x[264]^x[252]^x[251]^x[246]^x[245]^x[242]^x[240]^x[239]^x[236]^x[234]^x[231]^x[228]^x[225]^x[157]^x[156]^x[154]^x[146]^x[132]^x[92]^x[91]^x[82]^x[80]^x[79]^x[73]^x[71]^x[68]^x[67]^x[28];
	y[27]=x[307]^x[296]^x[285]^x[283]^x[263]^x[251]^x[250]^x[245]^x[244]^x[241]^x[239]^x[238]^x[235]^x[233]^x[230]^x[227]^x[224]^x[156]^x[155]^x[153]^x[145]^x[131]^x[91]^x[90]^x[81]^x[79]^x[78]^x[72]^x[70]^x[67]^x[66]^x[27];
	y[26]=x[372]^x[371]^x[361]^x[319]^x[318]^x[307]^x[284]^x[282]^x[262]^x[255]^x[250]^x[249]^x[244]^x[243]^x[240]^x[238]^x[237]^x[232]^x[229]^x[226]^x[155]^x[154]^x[152]^x[144]^x[130]^x[95]^x[90]^x[83]^x[80]^x[78]^x[74]^x[69]^x[68]^x[66]^x[53]^x[26];
	y[25]=x[371]^x[370]^x[360]^x[318]^x[317]^x[306]^x[283]^x[281]^x[261]^x[254]^x[249]^x[248]^x[243]^x[242]^x[239]^x[237]^x[236]^x[231]^x[228]^x[225]^x[154]^x[153]^x[151]^x[143]^x[129]^x[94]^x[89]^x[82]^x[79]^x[77]^x[73]^x[68]^x[67]^x[65]^x[63]^x[52]^x[42]^x[25];
	y[24]=x[370]^x[369]^x[359]^x[317]^x[316]^x[305]^x[282]^x[280]^x[260]^x[253]^x[248]^x[247]^x[242]^x[241]^x[238]^x[236]^x[235]^x[230]^x[227]^x[224]^x[153]^x[152]^x[150]^x[142]^x[128]^x[93]^x[88]^x[81]^x[78]^x[76]^x[72]^x[67]^x[66]^x[64]^x[62]^x[51]^x[41]^x[24];
	y[23]=x[369]^x[368]^x[358]^x[316]^x[315]^x[304]^x[303]^x[292]^x[281]^x[279]^x[259]^x[252]^x[247]^x[246]^x[241]^x[240]^x[237]^x[235]^x[229]^x[226]^x[152]^x[151]^x[141]^x[92]^x[87]^x[80]^x[77]^x[75]^x[74]^x[71]^x[68]^x[66]^x[65]^x[61]^x[50]^x[40]^x[23];
	y[22]=x[368]^x[367]^x[357]^x[315]^x[314]^x[303]^x[302]^x[291]^x[280]^x[278]^x[258]^x[251]^x[246]^x[245]^x[240]^x[239]^x[236]^x[234]^x[228]^x[225]^x[151]^x[150]^x[140]^x[91]^x[86]^x[79]^x[76]^x[74]^x[73]^x[70]^x[67]^x[65]^x[64]^x[60]^x[49]^x[39]^x[22];
	y[21]=x[373]^x[366]^x[362]^x[314]^x[313]^x[302]^x[301]^x[290]^x[279]^x[277]^x[257]^x[250]^x[245]^x[244]^x[239]^x[238]^x[235]^x[233]^x[227]^x[224]^x[213]^x[202]^x[150]^x[149]^x[139]^x[138]^x[90]^x[85]^x[78]^x[75]^x[73]^x[72]^x[69]^x[66]^x[64]^x[59]^x[48]^x[38]^x[21];
	y[20]=x[382]^x[376]^x[278]^x[276]^x[256]^x[255]^x[249]^x[244]^x[243]^x[238]^x[237]^x[232]^x[226]^x[222]^x[158]^x[149]^x[148]^x[146]^x[138]^x[137]^x[95]^x[84]^x[83]^x[72]^x[58]^x[37]^x[20];
	y[19]=x[381]^x[375]^x[287]^x[277]^x[275]^x[266]^x[254]^x[248]^x[243]^x[242]^x[237]^x[236]^x[231]^x[225]^x[221]^x[157]^x[148]^x[147]^x[145]^x[137]^x[136]^x[94]^x[83]^x[82]^x[71]^x[19];
	y[18]=x[380]^x[374]^x[286]^x[276]^x[274]^x[265]^x[253]^x[247]^x[242]^x[241]^x[236]^x[235]^x[230]^x[224]^x[220]^x[156]^x[147]^x[146]^x[144]^x[136]^x[135]^x[93]^x[82]^x[81]^x[70]^x[18];
	y[17]=x[379]^x[373]^x[363]^x[362]^x[352]^x[309]^x[298]^x[285]^x[275]^x[273]^x[264]^x[252]^x[246]^x[241]^x[240]^x[235]^x[229]^x[219]^x[155]^x[146]^x[145]^x[143]^x[135]^x[134]^x[92]^x[81]^x[80]^x[74]^x[69]^x[68]^x[17];
	y[16]=x[378]^x[372]^x[361]^x[308]^x[297]^x[284]^x[274]^x[272]^x[263]^x[251]^x[245]^x[240]^x[239]^x[234]^x[228]^x[218]^x[154]^x[145]^x[144]^x[142]^x[134]^x[133]^x[91]^x[80]^x[79]^x[73]^x[68]^x[67]^x[16];
	y[15]=x[377]^x[371]^x[360]^x[307]^x[296]^x[283]^x[273]^x[271]^x[262]^x[250]^x[244]^x[239]^x[238]^x[233]^x[227]^x[217]^x[153]^x[144]^x[143]^x[141]^x[133]^x[132]^x[90]^x[79]^x[78]^x[72]^x[67]^x[66]^x[42]^x[15];
	y[14]=x[376]^x[370]^x[359]^x[306]^x[295]^x[282]^x[272]^x[270]^x[261]^x[249]^x[243]^x[238]^x[237]^x[232]^x[226]^x[216]^x[152]^x[143]^x[142]^x[140]^x[132]^x[131]^x[89]^x[78]^x[77]^x[71]^x[66]^x[65]^x[41]^x[14];
	y[13]=x[375]^x[369]^x[358]^x[305]^x[294]^x[281]^x[271]^x[269]^x[260]^x[248]^x[242]^x[237]^x[236]^x[231]^x[225]^x[215]^x[151]^x[142]^x[141]^x[139]^x[131]^x[130]^x[88]^x[77]^x[76]^x[70]^x[65]^x[64]^x[40]^x[13];
	y[12]=x[374]^x[368]^x[357]^x[304]^x[293]^x[280]^x[270]^x[268]^x[259]^x[247]^x[241]^x[236]^x[235]^x[230]^x[224]^x[214]^x[150]^x[141]^x[140]^x[130]^x[129]^x[87]^x[76]^x[75]^x[69]^x[64]^x[39]^x[12];
	y[11]=x[363]^x[352]^x[279]^x[269]^x[267]^x[258]^x[246]^x[240]^x[235]^x[229]^x[203]^x[192]^x[140]^x[139]^x[129]^x[128]^x[86]^x[75]^x[38]^x[11];
	y[10]=x[278]^x[268]^x[266]^x[257]^x[245]^x[239]^x[234]^x[228]^x[139]^x[138]^x[128]^x[85]^x[74]^x[37]^x[10];
	y[9]=x[382]^x[376]^x[371]^x[365]^x[277]^x[267]^x[265]^x[256]^x[244]^x[238]^x[233]^x[227]^x[222]^x[211]^x[159]^x[147]^x[137]^x[135]^x[84]^x[73]^x[9];
	y[8]=x[381]^x[375]^x[370]^x[364]^x[287]^x[276]^x[264]^x[243]^x[237]^x[232]^x[226]^x[221]^x[210]^x[158]^x[146]^x[136]^x[134]^x[83]^x[72]^x[8];
	y[7]=x[380]^x[374]^x[369]^x[363]^x[286]^x[275]^x[263]^x[242]^x[236]^x[231]^x[225]^x[220]^x[209]^x[157]^x[145]^x[135]^x[133]^x[82]^x[71]^x[7];
	y[6]=x[379]^x[373]^x[368]^x[362]^x[285]^x[274]^x[262]^x[241]^x[235]^x[230]^x[224]^x[219]^x[208]^x[156]^x[144]^x[134]^x[132]^x[81]^x[70]^x[6];
	y[5]=x[378]^x[372]^x[367]^x[361]^x[309]^x[298]^x[284]^x[273]^x[261]^x[240]^x[229]^x[218]^x[207]^x[155]^x[143]^x[133]^x[131]^x[80]^x[74]^x[69]^x[68]^x[43]^x[32]^x[5];
	y[4]=x[377]^x[371]^x[366]^x[360]^x[308]^x[297]^x[283]^x[272]^x[260]^x[239]^x[228]^x[217]^x[206]^x[154]^x[142]^x[132]^x[130]^x[79]^x[73]^x[68]^x[67]^x[42]^x[4];
	y[3]=x[376]^x[370]^x[365]^x[359]^x[307]^x[296]^x[282]^x[271]^x[259]^x[238]^x[227]^x[216]^x[205]^x[153]^x[141]^x[131]^x[129]^x[78]^x[72]^x[67]^x[66]^x[41]^x[3];
	y[2]=x[375]^x[369]^x[364]^x[358]^x[306]^x[295]^x[281]^x[270]^x[258]^x[237]^x[226]^x[215]^x[204]^x[152]^x[140]^x[130]^x[128]^x[77]^x[71]^x[66]^x[65]^x[40]^x[2];
	y[1]=x[374]^x[368]^x[363]^x[357]^x[305]^x[294]^x[280]^x[269]^x[257]^x[236]^x[225]^x[214]^x[203]^x[151]^x[139]^x[129]^x[76]^x[70]^x[65]^x[64]^x[39]^x[1];
	y[0]=x[304]^x[293]^x[279]^x[268]^x[256]^x[235]^x[224]^x[150]^x[128]^x[75]^x[69]^x[64]^x[38]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint40(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[373]^x[362]^x[351]^x[345]^x[340]^x[334]^x[255]^x[236]^x[235]^x[225]^x[223]^x[222]^x[217]^x[216]^x[213]^x[211]^x[210]^x[207]^x[205]^x[204]^x[202]^x[199]^x[196]^x[193]^x[191]^x[180]^x[159]^x[153]^x[127]^x[125]^x[117]^x[116]^x[107]^x[104]^x[103]^x[96]^x[63]^x[62]^x[53]^x[51]^x[50]^x[42]^x[39]^x[26];
	y[30]=x[382]^x[372]^x[361]^x[254]^x[235]^x[234]^x[224]^x[222]^x[221]^x[216]^x[215]^x[212]^x[210]^x[209]^x[206]^x[204]^x[203]^x[201]^x[198]^x[195]^x[192]^x[158]^x[152]^x[127]^x[126]^x[124]^x[116]^x[102]^x[62]^x[61]^x[52]^x[50]^x[49]^x[41]^x[38];
	y[29]=x[381]^x[371]^x[360]^x[277]^x[266]^x[255]^x[253]^x[233]^x[221]^x[220]^x[215]^x[214]^x[211]^x[209]^x[208]^x[205]^x[203]^x[200]^x[197]^x[194]^x[157]^x[151]^x[126]^x[125]^x[123]^x[115]^x[101]^x[61]^x[60]^x[51]^x[49]^x[48]^x[42]^x[40]^x[37]^x[36];
	y[28]=x[380]^x[370]^x[359]^x[276]^x[265]^x[254]^x[252]^x[232]^x[220]^x[219]^x[214]^x[213]^x[210]^x[208]^x[207]^x[204]^x[202]^x[199]^x[196]^x[193]^x[156]^x[150]^x[125]^x[124]^x[122]^x[114]^x[100]^x[60]^x[59]^x[50]^x[48]^x[47]^x[41]^x[39]^x[36]^x[35];
	y[27]=x[379]^x[369]^x[358]^x[275]^x[264]^x[253]^x[251]^x[231]^x[219]^x[218]^x[213]^x[212]^x[209]^x[207]^x[206]^x[203]^x[201]^x[198]^x[195]^x[192]^x[155]^x[149]^x[124]^x[123]^x[121]^x[113]^x[99]^x[59]^x[58]^x[49]^x[47]^x[46]^x[40]^x[38]^x[35]^x[34];
	y[26]=x[378]^x[368]^x[357]^x[340]^x[339]^x[329]^x[287]^x[286]^x[275]^x[252]^x[250]^x[230]^x[223]^x[218]^x[217]^x[212]^x[211]^x[208]^x[206]^x[205]^x[200]^x[197]^x[194]^x[154]^x[148]^x[123]^x[122]^x[120]^x[112]^x[98]^x[63]^x[58]^x[51]^x[48]^x[46]^x[42]^x[37]^x[36]^x[34]^x[21];
	y[25]=x[377]^x[367]^x[356]^x[339]^x[338]^x[328]^x[286]^x[285]^x[274]^x[251]^x[249]^x[229]^x[222]^x[217]^x[216]^x[211]^x[210]^x[207]^x[205]^x[204]^x[199]^x[196]^x[193]^x[153]^x[147]^x[122]^x[121]^x[119]^x[111]^x[97]^x[62]^x[57]^x[50]^x[47]^x[45]^x[41]^x[36]^x[35]^x[33]^x[31]^x[20]^x[10];
	y[24]=x[376]^x[366]^x[355]^x[338]^x[337]^x[327]^x[285]^x[284]^x[273]^x[250]^x[248]^x[228]^x[221]^x[216]^x[215]^x[210]^x[209]^x[206]^x[204]^x[203]^x[198]^x[195]^x[192]^x[152]^x[146]^x[121]^x[120]^x[118]^x[110]^x[96]^x[61]^x[56]^x[49]^x[46]^x[44]^x[40]^x[35]^x[34]^x[32]^x[30]^x[19]^x[9];
	y[23]=x[375]^x[365]^x[354]^x[337]^x[336]^x[326]^x[284]^x[283]^x[272]^x[271]^x[260]^x[249]^x[247]^x[227]^x[220]^x[215]^x[214]^x[209]^x[208]^x[205]^x[203]^x[197]^x[194]^x[151]^x[145]^x[120]^x[119]^x[109]^x[60]^x[55]^x[48]^x[45]^x[43]^x[42]^x[39]^x[36]^x[34]^x[33]^x[29]^x[18]^x[8];
	y[22]=x[374]^x[364]^x[353]^x[336]^x[335]^x[325]^x[283]^x[282]^x[271]^x[270]^x[259]^x[248]^x[246]^x[226]^x[219]^x[214]^x[213]^x[208]^x[207]^x[204]^x[202]^x[196]^x[193]^x[150]^x[144]^x[119]^x[118]^x[108]^x[59]^x[54]^x[47]^x[44]^x[42]^x[41]^x[38]^x[35]^x[33]^x[32]^x[28]^x[17]^x[7];
	y[21]=x[373]^x[363]^x[352]^x[341]^x[334]^x[330]^x[282]^x[281]^x[270]^x[269]^x[258]^x[247]^x[245]^x[225]^x[218]^x[213]^x[212]^x[207]^x[206]^x[203]^x[201]^x[195]^x[192]^x[181]^x[170]^x[149]^x[143]^x[118]^x[117]^x[107]^x[106]^x[58]^x[53]^x[46]^x[43]^x[41]^x[40]^x[37]^x[34]^x[32]^x[27]^x[16]^x[6];
	y[20]=x[383]^x[372]^x[350]^x[344]^x[246]^x[244]^x[224]^x[223]^x[217]^x[212]^x[211]^x[206]^x[205]^x[200]^x[194]^x[190]^x[148]^x[142]^x[126]^x[117]^x[116]^x[114]^x[106]^x[105]^x[63]^x[52]^x[51]^x[40]^x[26]^x[5];
	y[19]=x[382]^x[371]^x[349]^x[343]^x[255]^x[245]^x[243]^x[234]^x[222]^x[216]^x[211]^x[210]^x[205]^x[204]^x[199]^x[193]^x[189]^x[147]^x[141]^x[125]^x[116]^x[115]^x[113]^x[105]^x[104]^x[62]^x[51]^x[50]^x[39];
	y[18]=x[381]^x[370]^x[348]^x[342]^x[254]^x[244]^x[242]^x[233]^x[221]^x[215]^x[210]^x[209]^x[204]^x[203]^x[198]^x[192]^x[188]^x[146]^x[140]^x[124]^x[115]^x[114]^x[112]^x[104]^x[103]^x[61]^x[50]^x[49]^x[38];
	y[17]=x[380]^x[369]^x[347]^x[341]^x[331]^x[330]^x[320]^x[277]^x[266]^x[253]^x[243]^x[241]^x[232]^x[220]^x[214]^x[209]^x[208]^x[203]^x[197]^x[187]^x[145]^x[139]^x[123]^x[114]^x[113]^x[111]^x[103]^x[102]^x[60]^x[49]^x[48]^x[42]^x[37]^x[36];
	y[16]=x[379]^x[368]^x[346]^x[340]^x[329]^x[276]^x[265]^x[252]^x[242]^x[240]^x[231]^x[219]^x[213]^x[208]^x[207]^x[202]^x[196]^x[186]^x[144]^x[138]^x[122]^x[113]^x[112]^x[110]^x[102]^x[101]^x[59]^x[48]^x[47]^x[41]^x[36]^x[35];
	y[15]=x[378]^x[367]^x[345]^x[339]^x[328]^x[275]^x[264]^x[251]^x[241]^x[239]^x[230]^x[218]^x[212]^x[207]^x[206]^x[201]^x[195]^x[185]^x[143]^x[137]^x[121]^x[112]^x[111]^x[109]^x[101]^x[100]^x[58]^x[47]^x[46]^x[40]^x[35]^x[34]^x[10];
	y[14]=x[377]^x[366]^x[344]^x[338]^x[327]^x[274]^x[263]^x[250]^x[240]^x[238]^x[229]^x[217]^x[211]^x[206]^x[205]^x[200]^x[194]^x[184]^x[142]^x[136]^x[120]^x[111]^x[110]^x[108]^x[100]^x[99]^x[57]^x[46]^x[45]^x[39]^x[34]^x[33]^x[9];
	y[13]=x[376]^x[365]^x[343]^x[337]^x[326]^x[273]^x[262]^x[249]^x[239]^x[237]^x[228]^x[216]^x[210]^x[205]^x[204]^x[199]^x[193]^x[183]^x[141]^x[135]^x[119]^x[110]^x[109]^x[107]^x[99]^x[98]^x[56]^x[45]^x[44]^x[38]^x[33]^x[32]^x[8];
	y[12]=x[375]^x[364]^x[342]^x[336]^x[325]^x[272]^x[261]^x[248]^x[238]^x[236]^x[227]^x[215]^x[209]^x[204]^x[203]^x[198]^x[192]^x[182]^x[140]^x[134]^x[118]^x[109]^x[108]^x[98]^x[97]^x[55]^x[44]^x[43]^x[37]^x[32]^x[7];
	y[11]=x[374]^x[363]^x[331]^x[320]^x[247]^x[237]^x[235]^x[226]^x[214]^x[208]^x[203]^x[197]^x[171]^x[160]^x[139]^x[133]^x[108]^x[107]^x[97]^x[96]^x[54]^x[43]^x[6];
	y[10]=x[373]^x[362]^x[246]^x[236]^x[234]^x[225]^x[213]^x[207]^x[202]^x[196]^x[138]^x[132]^x[107]^x[106]^x[96]^x[53]^x[42]^x[5];
	y[9]=x[372]^x[361]^x[350]^x[344]^x[339]^x[333]^x[245]^x[235]^x[233]^x[224]^x[212]^x[206]^x[201]^x[195]^x[190]^x[179]^x[137]^x[131]^x[127]^x[115]^x[105]^x[103]^x[52]^x[41];
	y[8]=x[371]^x[360]^x[349]^x[343]^x[338]^x[332]^x[255]^x[244]^x[232]^x[211]^x[205]^x[200]^x[194]^x[189]^x[178]^x[136]^x[130]^x[126]^x[114]^x[104]^x[102]^x[51]^x[40];
	y[7]=x[370]^x[359]^x[348]^x[342]^x[337]^x[331]^x[254]^x[243]^x[231]^x[210]^x[204]^x[199]^x[193]^x[188]^x[177]^x[135]^x[129]^x[125]^x[113]^x[103]^x[101]^x[50]^x[39];
	y[6]=x[369]^x[358]^x[347]^x[341]^x[336]^x[330]^x[253]^x[242]^x[230]^x[209]^x[203]^x[198]^x[192]^x[187]^x[176]^x[134]^x[128]^x[124]^x[112]^x[102]^x[100]^x[49]^x[38];
	y[5]=x[368]^x[357]^x[346]^x[340]^x[335]^x[329]^x[277]^x[266]^x[252]^x[241]^x[229]^x[208]^x[197]^x[186]^x[175]^x[133]^x[123]^x[111]^x[101]^x[99]^x[48]^x[42]^x[37]^x[36]^x[11]^x[0];
	y[4]=x[367]^x[356]^x[345]^x[339]^x[334]^x[328]^x[276]^x[265]^x[251]^x[240]^x[228]^x[207]^x[196]^x[185]^x[174]^x[132]^x[122]^x[110]^x[100]^x[98]^x[47]^x[41]^x[36]^x[35]^x[10];
	y[3]=x[366]^x[355]^x[344]^x[338]^x[333]^x[327]^x[275]^x[264]^x[250]^x[239]^x[227]^x[206]^x[195]^x[184]^x[173]^x[131]^x[121]^x[109]^x[99]^x[97]^x[46]^x[40]^x[35]^x[34]^x[9];
	y[2]=x[365]^x[354]^x[343]^x[337]^x[332]^x[326]^x[274]^x[263]^x[249]^x[238]^x[226]^x[205]^x[194]^x[183]^x[172]^x[130]^x[120]^x[108]^x[98]^x[96]^x[45]^x[39]^x[34]^x[33]^x[8];
	y[1]=x[364]^x[353]^x[342]^x[336]^x[331]^x[325]^x[273]^x[262]^x[248]^x[237]^x[225]^x[204]^x[193]^x[182]^x[171]^x[129]^x[119]^x[107]^x[97]^x[44]^x[38]^x[33]^x[32]^x[7];
	y[0]=x[363]^x[352]^x[272]^x[261]^x[247]^x[236]^x[224]^x[203]^x[192]^x[128]^x[118]^x[96]^x[43]^x[37]^x[32]^x[6];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint41(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[378]^x[368]^x[357]^x[351]^x[341]^x[330]^x[319]^x[313]^x[308]^x[302]^x[223]^x[204]^x[203]^x[193]^x[191]^x[190]^x[185]^x[184]^x[181]^x[179]^x[178]^x[175]^x[173]^x[172]^x[170]^x[167]^x[164]^x[161]^x[159]^x[154]^x[127]^x[121]^x[95]^x[93]^x[85]^x[84]^x[75]^x[72]^x[71]^x[64]^x[31]^x[30]^x[21]^x[19]^x[18]^x[10]^x[7];
	y[30]=x[350]^x[340]^x[329]^x[222]^x[203]^x[202]^x[192]^x[190]^x[189]^x[184]^x[183]^x[180]^x[178]^x[177]^x[174]^x[172]^x[171]^x[169]^x[166]^x[163]^x[160]^x[126]^x[120]^x[95]^x[94]^x[92]^x[84]^x[70]^x[30]^x[29]^x[20]^x[18]^x[17]^x[9]^x[6];
	y[29]=x[349]^x[339]^x[328]^x[245]^x[234]^x[223]^x[221]^x[201]^x[189]^x[188]^x[183]^x[182]^x[179]^x[177]^x[176]^x[173]^x[171]^x[168]^x[165]^x[162]^x[125]^x[119]^x[94]^x[93]^x[91]^x[83]^x[69]^x[29]^x[28]^x[19]^x[17]^x[16]^x[10]^x[8]^x[5]^x[4];
	y[28]=x[348]^x[338]^x[327]^x[244]^x[233]^x[222]^x[220]^x[200]^x[188]^x[187]^x[182]^x[181]^x[178]^x[176]^x[175]^x[172]^x[170]^x[167]^x[164]^x[161]^x[124]^x[118]^x[93]^x[92]^x[90]^x[82]^x[68]^x[28]^x[27]^x[18]^x[16]^x[15]^x[9]^x[7]^x[4]^x[3];
	y[27]=x[347]^x[337]^x[326]^x[243]^x[232]^x[221]^x[219]^x[199]^x[187]^x[186]^x[181]^x[180]^x[177]^x[175]^x[174]^x[171]^x[169]^x[166]^x[163]^x[160]^x[123]^x[117]^x[92]^x[91]^x[89]^x[81]^x[67]^x[27]^x[26]^x[17]^x[15]^x[14]^x[8]^x[6]^x[3]^x[2];
	y[26]=x[373]^x[363]^x[352]^x[346]^x[336]^x[325]^x[308]^x[307]^x[297]^x[255]^x[254]^x[243]^x[220]^x[218]^x[198]^x[191]^x[186]^x[185]^x[180]^x[179]^x[176]^x[174]^x[173]^x[168]^x[165]^x[162]^x[149]^x[143]^x[122]^x[116]^x[91]^x[90]^x[88]^x[80]^x[66]^x[31]^x[26]^x[19]^x[16]^x[14]^x[10]^x[5]^x[4]^x[2];
	y[25]=x[372]^x[345]^x[335]^x[324]^x[307]^x[306]^x[296]^x[254]^x[253]^x[242]^x[219]^x[217]^x[197]^x[190]^x[185]^x[184]^x[179]^x[178]^x[175]^x[173]^x[172]^x[167]^x[164]^x[161]^x[159]^x[153]^x[148]^x[142]^x[138]^x[132]^x[121]^x[115]^x[90]^x[89]^x[87]^x[79]^x[65]^x[30]^x[25]^x[18]^x[15]^x[13]^x[9]^x[4]^x[3]^x[1];
	y[24]=x[371]^x[344]^x[334]^x[323]^x[306]^x[305]^x[295]^x[253]^x[252]^x[241]^x[218]^x[216]^x[196]^x[189]^x[184]^x[183]^x[178]^x[177]^x[174]^x[172]^x[171]^x[166]^x[163]^x[160]^x[158]^x[152]^x[147]^x[141]^x[137]^x[131]^x[120]^x[114]^x[89]^x[88]^x[86]^x[78]^x[64]^x[29]^x[24]^x[17]^x[14]^x[12]^x[8]^x[3]^x[2]^x[0];
	y[23]=x[370]^x[343]^x[333]^x[322]^x[305]^x[304]^x[294]^x[252]^x[251]^x[240]^x[239]^x[228]^x[217]^x[215]^x[195]^x[188]^x[183]^x[182]^x[177]^x[176]^x[173]^x[171]^x[165]^x[162]^x[157]^x[151]^x[146]^x[140]^x[136]^x[130]^x[119]^x[113]^x[88]^x[87]^x[77]^x[28]^x[23]^x[16]^x[13]^x[11]^x[10]^x[7]^x[4]^x[2]^x[1];
	y[22]=x[369]^x[342]^x[332]^x[321]^x[304]^x[303]^x[293]^x[251]^x[250]^x[239]^x[238]^x[227]^x[216]^x[214]^x[194]^x[187]^x[182]^x[181]^x[176]^x[175]^x[172]^x[170]^x[164]^x[161]^x[156]^x[150]^x[145]^x[139]^x[135]^x[129]^x[118]^x[112]^x[87]^x[86]^x[76]^x[27]^x[22]^x[15]^x[12]^x[10]^x[9]^x[6]^x[3]^x[1]^x[0];
	y[21]=x[368]^x[341]^x[331]^x[320]^x[309]^x[302]^x[298]^x[250]^x[249]^x[238]^x[237]^x[226]^x[215]^x[213]^x[193]^x[186]^x[181]^x[180]^x[175]^x[174]^x[171]^x[169]^x[163]^x[160]^x[155]^x[144]^x[134]^x[128]^x[117]^x[111]^x[86]^x[85]^x[75]^x[74]^x[26]^x[21]^x[14]^x[11]^x[9]^x[8]^x[5]^x[2]^x[0];
	y[20]=x[378]^x[351]^x[340]^x[318]^x[312]^x[214]^x[212]^x[192]^x[191]^x[185]^x[180]^x[179]^x[174]^x[173]^x[168]^x[162]^x[158]^x[154]^x[148]^x[133]^x[116]^x[110]^x[94]^x[85]^x[84]^x[82]^x[74]^x[73]^x[31]^x[20]^x[19]^x[8];
	y[19]=x[350]^x[339]^x[317]^x[311]^x[223]^x[213]^x[211]^x[202]^x[190]^x[184]^x[179]^x[178]^x[173]^x[172]^x[167]^x[161]^x[157]^x[115]^x[109]^x[93]^x[84]^x[83]^x[81]^x[73]^x[72]^x[30]^x[19]^x[18]^x[7];
	y[18]=x[349]^x[338]^x[316]^x[310]^x[222]^x[212]^x[210]^x[201]^x[189]^x[183]^x[178]^x[177]^x[172]^x[171]^x[166]^x[160]^x[156]^x[114]^x[108]^x[92]^x[83]^x[82]^x[80]^x[72]^x[71]^x[29]^x[18]^x[17]^x[6];
	y[17]=x[348]^x[337]^x[315]^x[309]^x[299]^x[298]^x[288]^x[245]^x[234]^x[221]^x[211]^x[209]^x[200]^x[188]^x[182]^x[177]^x[176]^x[171]^x[165]^x[155]^x[113]^x[107]^x[91]^x[82]^x[81]^x[79]^x[71]^x[70]^x[28]^x[17]^x[16]^x[10]^x[5]^x[4];
	y[16]=x[347]^x[336]^x[314]^x[308]^x[297]^x[244]^x[233]^x[220]^x[210]^x[208]^x[199]^x[187]^x[181]^x[176]^x[175]^x[170]^x[164]^x[154]^x[112]^x[106]^x[90]^x[81]^x[80]^x[78]^x[70]^x[69]^x[27]^x[16]^x[15]^x[9]^x[4]^x[3];
	y[15]=x[373]^x[362]^x[346]^x[335]^x[313]^x[307]^x[296]^x[243]^x[232]^x[219]^x[209]^x[207]^x[198]^x[186]^x[180]^x[175]^x[174]^x[169]^x[163]^x[153]^x[138]^x[132]^x[111]^x[105]^x[89]^x[80]^x[79]^x[77]^x[69]^x[68]^x[26]^x[15]^x[14]^x[8]^x[3]^x[2];
	y[14]=x[372]^x[361]^x[345]^x[334]^x[312]^x[306]^x[295]^x[242]^x[231]^x[218]^x[208]^x[206]^x[197]^x[185]^x[179]^x[174]^x[173]^x[168]^x[162]^x[152]^x[137]^x[131]^x[110]^x[104]^x[88]^x[79]^x[78]^x[76]^x[68]^x[67]^x[25]^x[14]^x[13]^x[7]^x[2]^x[1];
	y[13]=x[371]^x[360]^x[344]^x[333]^x[311]^x[305]^x[294]^x[241]^x[230]^x[217]^x[207]^x[205]^x[196]^x[184]^x[178]^x[173]^x[172]^x[167]^x[161]^x[151]^x[136]^x[130]^x[109]^x[103]^x[87]^x[78]^x[77]^x[75]^x[67]^x[66]^x[24]^x[13]^x[12]^x[6]^x[1]^x[0];
	y[12]=x[370]^x[359]^x[343]^x[332]^x[310]^x[304]^x[293]^x[240]^x[229]^x[216]^x[206]^x[204]^x[195]^x[183]^x[177]^x[172]^x[171]^x[166]^x[160]^x[150]^x[135]^x[129]^x[108]^x[102]^x[86]^x[77]^x[76]^x[66]^x[65]^x[23]^x[12]^x[11]^x[5]^x[0];
	y[11]=x[369]^x[358]^x[342]^x[331]^x[299]^x[288]^x[215]^x[205]^x[203]^x[194]^x[182]^x[176]^x[171]^x[165]^x[139]^x[134]^x[107]^x[101]^x[76]^x[75]^x[65]^x[64]^x[22]^x[11];
	y[10]=x[368]^x[357]^x[341]^x[330]^x[214]^x[204]^x[202]^x[193]^x[181]^x[175]^x[170]^x[164]^x[133]^x[106]^x[100]^x[75]^x[74]^x[64]^x[21]^x[10];
	y[9]=x[340]^x[329]^x[318]^x[312]^x[307]^x[301]^x[213]^x[203]^x[201]^x[192]^x[180]^x[174]^x[169]^x[163]^x[158]^x[147]^x[105]^x[99]^x[95]^x[83]^x[73]^x[71]^x[20]^x[9];
	y[8]=x[339]^x[328]^x[317]^x[311]^x[306]^x[300]^x[223]^x[212]^x[200]^x[179]^x[173]^x[168]^x[162]^x[157]^x[146]^x[104]^x[98]^x[94]^x[82]^x[72]^x[70]^x[19]^x[8];
	y[7]=x[338]^x[327]^x[316]^x[310]^x[305]^x[299]^x[222]^x[211]^x[199]^x[178]^x[172]^x[167]^x[161]^x[156]^x[145]^x[103]^x[97]^x[93]^x[81]^x[71]^x[69]^x[18]^x[7];
	y[6]=x[337]^x[326]^x[315]^x[309]^x[304]^x[298]^x[221]^x[210]^x[198]^x[177]^x[171]^x[166]^x[160]^x[155]^x[144]^x[102]^x[96]^x[92]^x[80]^x[70]^x[68]^x[17]^x[6];
	y[5]=x[374]^x[352]^x[336]^x[325]^x[314]^x[308]^x[303]^x[297]^x[245]^x[234]^x[220]^x[209]^x[197]^x[176]^x[165]^x[154]^x[143]^x[139]^x[133]^x[128]^x[101]^x[91]^x[79]^x[69]^x[67]^x[16]^x[10]^x[5]^x[4];
	y[4]=x[373]^x[362]^x[335]^x[324]^x[313]^x[307]^x[302]^x[296]^x[244]^x[233]^x[219]^x[208]^x[196]^x[175]^x[164]^x[153]^x[142]^x[138]^x[132]^x[100]^x[90]^x[78]^x[68]^x[66]^x[15]^x[9]^x[4]^x[3];
	y[3]=x[372]^x[361]^x[334]^x[323]^x[312]^x[306]^x[301]^x[295]^x[243]^x[232]^x[218]^x[207]^x[195]^x[174]^x[163]^x[152]^x[141]^x[137]^x[131]^x[99]^x[89]^x[77]^x[67]^x[65]^x[14]^x[8]^x[3]^x[2];
	y[2]=x[371]^x[360]^x[333]^x[322]^x[311]^x[305]^x[300]^x[294]^x[242]^x[231]^x[217]^x[206]^x[194]^x[173]^x[162]^x[151]^x[140]^x[136]^x[130]^x[98]^x[88]^x[76]^x[66]^x[64]^x[13]^x[7]^x[2]^x[1];
	y[1]=x[370]^x[359]^x[332]^x[321]^x[310]^x[304]^x[299]^x[293]^x[241]^x[230]^x[216]^x[205]^x[193]^x[172]^x[161]^x[150]^x[139]^x[135]^x[129]^x[97]^x[87]^x[75]^x[65]^x[12]^x[6]^x[1]^x[0];
	y[0]=x[369]^x[358]^x[331]^x[320]^x[240]^x[229]^x[215]^x[204]^x[192]^x[171]^x[160]^x[134]^x[128]^x[96]^x[86]^x[64]^x[11]^x[5]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint42(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[381]^x[373]^x[372]^x[371]^x[363]^x[361]^x[359]^x[352]^x[346]^x[336]^x[325]^x[319]^x[309]^x[298]^x[287]^x[281]^x[276]^x[270]^x[191]^x[172]^x[171]^x[161]^x[127]^x[122]^x[95]^x[89]^x[63]^x[61]^x[53]^x[52]^x[43]^x[40]^x[39]^x[32];
	y[30]=x[383]^x[382]^x[380]^x[372]^x[371]^x[370]^x[360]^x[358]^x[318]^x[308]^x[297]^x[190]^x[171]^x[170]^x[160]^x[94]^x[88]^x[63]^x[62]^x[60]^x[52]^x[38];
	y[29]=x[382]^x[381]^x[379]^x[373]^x[371]^x[370]^x[369]^x[367]^x[362]^x[359]^x[357]^x[356]^x[317]^x[307]^x[296]^x[213]^x[202]^x[191]^x[189]^x[169]^x[93]^x[87]^x[62]^x[61]^x[59]^x[51]^x[37];
	y[28]=x[381]^x[380]^x[378]^x[372]^x[370]^x[369]^x[368]^x[366]^x[361]^x[358]^x[356]^x[355]^x[316]^x[306]^x[295]^x[212]^x[201]^x[190]^x[188]^x[168]^x[92]^x[86]^x[61]^x[60]^x[58]^x[50]^x[36];
	y[27]=x[380]^x[379]^x[377]^x[371]^x[369]^x[368]^x[367]^x[365]^x[360]^x[357]^x[355]^x[354]^x[315]^x[305]^x[294]^x[211]^x[200]^x[189]^x[187]^x[167]^x[91]^x[85]^x[60]^x[59]^x[57]^x[49]^x[35];
	y[26]=x[383]^x[382]^x[379]^x[378]^x[377]^x[371]^x[368]^x[367]^x[366]^x[365]^x[356]^x[354]^x[341]^x[331]^x[320]^x[314]^x[304]^x[293]^x[276]^x[275]^x[265]^x[223]^x[222]^x[211]^x[188]^x[186]^x[166]^x[117]^x[111]^x[90]^x[84]^x[59]^x[58]^x[56]^x[48]^x[34];
	y[25]=x[382]^x[381]^x[378]^x[377]^x[376]^x[370]^x[367]^x[366]^x[365]^x[364]^x[355]^x[353]^x[340]^x[313]^x[303]^x[292]^x[275]^x[274]^x[264]^x[222]^x[221]^x[210]^x[187]^x[185]^x[165]^x[127]^x[121]^x[116]^x[110]^x[106]^x[100]^x[89]^x[83]^x[58]^x[57]^x[55]^x[47]^x[33];
	y[24]=x[381]^x[380]^x[377]^x[376]^x[375]^x[369]^x[366]^x[365]^x[364]^x[363]^x[354]^x[352]^x[339]^x[312]^x[302]^x[291]^x[274]^x[273]^x[263]^x[221]^x[220]^x[209]^x[186]^x[184]^x[164]^x[126]^x[120]^x[115]^x[109]^x[105]^x[99]^x[88]^x[82]^x[57]^x[56]^x[54]^x[46]^x[32];
	y[23]=x[380]^x[379]^x[376]^x[375]^x[374]^x[373]^x[368]^x[367]^x[365]^x[364]^x[363]^x[362]^x[356]^x[353]^x[338]^x[311]^x[301]^x[290]^x[273]^x[272]^x[262]^x[220]^x[219]^x[208]^x[207]^x[196]^x[185]^x[183]^x[163]^x[125]^x[119]^x[114]^x[108]^x[104]^x[98]^x[87]^x[81]^x[56]^x[55]^x[45];
	y[22]=x[379]^x[378]^x[375]^x[374]^x[373]^x[372]^x[367]^x[366]^x[364]^x[363]^x[362]^x[361]^x[355]^x[352]^x[337]^x[310]^x[300]^x[289]^x[272]^x[271]^x[261]^x[219]^x[218]^x[207]^x[206]^x[195]^x[184]^x[182]^x[162]^x[124]^x[118]^x[113]^x[107]^x[103]^x[97]^x[86]^x[80]^x[55]^x[54]^x[44];
	y[21]=x[378]^x[377]^x[374]^x[373]^x[372]^x[371]^x[366]^x[365]^x[363]^x[361]^x[360]^x[354]^x[336]^x[309]^x[299]^x[288]^x[277]^x[270]^x[266]^x[218]^x[217]^x[206]^x[205]^x[194]^x[183]^x[181]^x[161]^x[123]^x[112]^x[102]^x[96]^x[85]^x[79]^x[54]^x[53]^x[43]^x[42];
	y[20]=x[382]^x[373]^x[372]^x[362]^x[360]^x[346]^x[319]^x[308]^x[286]^x[280]^x[182]^x[180]^x[160]^x[126]^x[122]^x[116]^x[101]^x[84]^x[78]^x[62]^x[53]^x[52]^x[50]^x[42]^x[41];
	y[19]=x[381]^x[372]^x[371]^x[361]^x[359]^x[318]^x[307]^x[285]^x[279]^x[191]^x[181]^x[179]^x[170]^x[125]^x[83]^x[77]^x[61]^x[52]^x[51]^x[49]^x[41]^x[40];
	y[18]=x[380]^x[371]^x[370]^x[360]^x[358]^x[317]^x[306]^x[284]^x[278]^x[190]^x[180]^x[178]^x[169]^x[124]^x[82]^x[76]^x[60]^x[51]^x[50]^x[48]^x[40]^x[39];
	y[17]=x[379]^x[373]^x[370]^x[369]^x[367]^x[362]^x[359]^x[357]^x[356]^x[316]^x[305]^x[283]^x[277]^x[267]^x[266]^x[256]^x[213]^x[202]^x[189]^x[179]^x[177]^x[168]^x[123]^x[81]^x[75]^x[59]^x[50]^x[49]^x[47]^x[39]^x[38];
	y[16]=x[378]^x[372]^x[369]^x[368]^x[366]^x[361]^x[358]^x[356]^x[355]^x[315]^x[304]^x[282]^x[276]^x[265]^x[212]^x[201]^x[188]^x[178]^x[176]^x[167]^x[122]^x[80]^x[74]^x[58]^x[49]^x[48]^x[46]^x[38]^x[37];
	y[15]=x[377]^x[371]^x[368]^x[367]^x[365]^x[360]^x[357]^x[355]^x[354]^x[341]^x[330]^x[314]^x[303]^x[281]^x[275]^x[264]^x[211]^x[200]^x[187]^x[177]^x[175]^x[166]^x[121]^x[106]^x[100]^x[79]^x[73]^x[57]^x[48]^x[47]^x[45]^x[37]^x[36];
	y[14]=x[376]^x[370]^x[367]^x[366]^x[364]^x[359]^x[356]^x[354]^x[353]^x[340]^x[329]^x[313]^x[302]^x[280]^x[274]^x[263]^x[210]^x[199]^x[186]^x[176]^x[174]^x[165]^x[120]^x[105]^x[99]^x[78]^x[72]^x[56]^x[47]^x[46]^x[44]^x[36]^x[35];
	y[13]=x[375]^x[369]^x[366]^x[365]^x[363]^x[358]^x[355]^x[353]^x[352]^x[339]^x[328]^x[312]^x[301]^x[279]^x[273]^x[262]^x[209]^x[198]^x[185]^x[175]^x[173]^x[164]^x[119]^x[104]^x[98]^x[77]^x[71]^x[55]^x[46]^x[45]^x[43]^x[35]^x[34];
	y[12]=x[374]^x[368]^x[365]^x[364]^x[357]^x[354]^x[352]^x[338]^x[327]^x[311]^x[300]^x[278]^x[272]^x[261]^x[208]^x[197]^x[184]^x[174]^x[172]^x[163]^x[118]^x[103]^x[97]^x[76]^x[70]^x[54]^x[45]^x[44]^x[34]^x[33];
	y[11]=x[364]^x[363]^x[353]^x[337]^x[326]^x[310]^x[299]^x[267]^x[256]^x[183]^x[173]^x[171]^x[162]^x[107]^x[102]^x[75]^x[69]^x[44]^x[43]^x[33]^x[32];
	y[10]=x[363]^x[362]^x[352]^x[336]^x[325]^x[309]^x[298]^x[182]^x[172]^x[170]^x[161]^x[101]^x[74]^x[68]^x[43]^x[42]^x[32];
	y[9]=x[383]^x[361]^x[308]^x[297]^x[286]^x[280]^x[275]^x[269]^x[181]^x[171]^x[169]^x[160]^x[126]^x[115]^x[73]^x[67]^x[63]^x[51]^x[41]^x[39];
	y[8]=x[382]^x[360]^x[307]^x[296]^x[285]^x[279]^x[274]^x[268]^x[191]^x[180]^x[168]^x[125]^x[114]^x[72]^x[66]^x[62]^x[50]^x[40]^x[38];
	y[7]=x[381]^x[359]^x[306]^x[295]^x[284]^x[278]^x[273]^x[267]^x[190]^x[179]^x[167]^x[124]^x[113]^x[71]^x[65]^x[61]^x[49]^x[39]^x[37];
	y[6]=x[380]^x[358]^x[305]^x[294]^x[283]^x[277]^x[272]^x[266]^x[189]^x[178]^x[166]^x[123]^x[112]^x[70]^x[64]^x[60]^x[48]^x[38]^x[36];
	y[5]=x[379]^x[373]^x[367]^x[362]^x[357]^x[356]^x[342]^x[320]^x[304]^x[293]^x[282]^x[276]^x[271]^x[265]^x[213]^x[202]^x[188]^x[177]^x[165]^x[122]^x[111]^x[107]^x[101]^x[96]^x[69]^x[59]^x[47]^x[37]^x[35];
	y[4]=x[378]^x[372]^x[366]^x[361]^x[356]^x[355]^x[341]^x[330]^x[303]^x[292]^x[281]^x[275]^x[270]^x[264]^x[212]^x[201]^x[187]^x[176]^x[164]^x[121]^x[110]^x[106]^x[100]^x[68]^x[58]^x[46]^x[36]^x[34];
	y[3]=x[377]^x[371]^x[365]^x[360]^x[355]^x[354]^x[340]^x[329]^x[302]^x[291]^x[280]^x[274]^x[269]^x[263]^x[211]^x[200]^x[186]^x[175]^x[163]^x[120]^x[109]^x[105]^x[99]^x[67]^x[57]^x[45]^x[35]^x[33];
	y[2]=x[376]^x[370]^x[364]^x[359]^x[354]^x[353]^x[339]^x[328]^x[301]^x[290]^x[279]^x[273]^x[268]^x[262]^x[210]^x[199]^x[185]^x[174]^x[162]^x[119]^x[108]^x[104]^x[98]^x[66]^x[56]^x[44]^x[34]^x[32];
	y[1]=x[375]^x[369]^x[363]^x[358]^x[353]^x[352]^x[338]^x[327]^x[300]^x[289]^x[278]^x[272]^x[267]^x[261]^x[209]^x[198]^x[184]^x[173]^x[161]^x[118]^x[107]^x[103]^x[97]^x[65]^x[55]^x[43]^x[33];
	y[0]=x[374]^x[368]^x[357]^x[352]^x[337]^x[326]^x[299]^x[288]^x[208]^x[197]^x[183]^x[172]^x[160]^x[102]^x[96]^x[64]^x[54]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint43(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[349]^x[341]^x[340]^x[339]^x[331]^x[329]^x[327]^x[320]^x[314]^x[304]^x[293]^x[287]^x[277]^x[266]^x[255]^x[249]^x[244]^x[238]^x[159]^x[140]^x[139]^x[129]^x[95]^x[90]^x[63]^x[57]^x[31]^x[29]^x[21]^x[20]^x[11]^x[8]^x[7]^x[0];
	y[30]=x[351]^x[350]^x[348]^x[340]^x[339]^x[338]^x[328]^x[326]^x[286]^x[276]^x[265]^x[158]^x[139]^x[138]^x[128]^x[62]^x[56]^x[31]^x[30]^x[28]^x[20]^x[6];
	y[29]=x[350]^x[349]^x[347]^x[341]^x[339]^x[338]^x[337]^x[335]^x[330]^x[327]^x[325]^x[324]^x[285]^x[275]^x[264]^x[181]^x[170]^x[159]^x[157]^x[137]^x[61]^x[55]^x[30]^x[29]^x[27]^x[19]^x[5];
	y[28]=x[349]^x[348]^x[346]^x[340]^x[338]^x[337]^x[336]^x[334]^x[329]^x[326]^x[324]^x[323]^x[284]^x[274]^x[263]^x[180]^x[169]^x[158]^x[156]^x[136]^x[60]^x[54]^x[29]^x[28]^x[26]^x[18]^x[4];
	y[27]=x[348]^x[347]^x[345]^x[339]^x[337]^x[336]^x[335]^x[333]^x[328]^x[325]^x[323]^x[322]^x[283]^x[273]^x[262]^x[179]^x[168]^x[157]^x[155]^x[135]^x[59]^x[53]^x[28]^x[27]^x[25]^x[17]^x[3];
	y[26]=x[351]^x[350]^x[347]^x[346]^x[345]^x[339]^x[336]^x[335]^x[334]^x[333]^x[324]^x[322]^x[309]^x[299]^x[288]^x[282]^x[272]^x[261]^x[244]^x[243]^x[233]^x[191]^x[190]^x[179]^x[156]^x[154]^x[134]^x[85]^x[79]^x[58]^x[52]^x[27]^x[26]^x[24]^x[16]^x[2];
	y[25]=x[350]^x[349]^x[346]^x[345]^x[344]^x[338]^x[335]^x[334]^x[333]^x[332]^x[323]^x[321]^x[308]^x[281]^x[271]^x[260]^x[243]^x[242]^x[232]^x[190]^x[189]^x[178]^x[155]^x[153]^x[133]^x[95]^x[89]^x[84]^x[78]^x[74]^x[68]^x[57]^x[51]^x[26]^x[25]^x[23]^x[15]^x[1];
	y[24]=x[349]^x[348]^x[345]^x[344]^x[343]^x[337]^x[334]^x[333]^x[332]^x[331]^x[322]^x[320]^x[307]^x[280]^x[270]^x[259]^x[242]^x[241]^x[231]^x[189]^x[188]^x[177]^x[154]^x[152]^x[132]^x[94]^x[88]^x[83]^x[77]^x[73]^x[67]^x[56]^x[50]^x[25]^x[24]^x[22]^x[14]^x[0];
	y[23]=x[348]^x[347]^x[344]^x[343]^x[342]^x[341]^x[336]^x[335]^x[333]^x[332]^x[331]^x[330]^x[324]^x[321]^x[306]^x[279]^x[269]^x[258]^x[241]^x[240]^x[230]^x[188]^x[187]^x[176]^x[175]^x[164]^x[153]^x[151]^x[131]^x[93]^x[87]^x[82]^x[76]^x[72]^x[66]^x[55]^x[49]^x[24]^x[23]^x[13];
	y[22]=x[347]^x[346]^x[343]^x[342]^x[341]^x[340]^x[335]^x[334]^x[332]^x[331]^x[330]^x[329]^x[323]^x[320]^x[305]^x[278]^x[268]^x[257]^x[240]^x[239]^x[229]^x[187]^x[186]^x[175]^x[174]^x[163]^x[152]^x[150]^x[130]^x[92]^x[86]^x[81]^x[75]^x[71]^x[65]^x[54]^x[48]^x[23]^x[22]^x[12];
	y[21]=x[346]^x[345]^x[342]^x[341]^x[340]^x[339]^x[334]^x[333]^x[331]^x[329]^x[328]^x[322]^x[304]^x[277]^x[267]^x[256]^x[245]^x[238]^x[234]^x[186]^x[185]^x[174]^x[173]^x[162]^x[151]^x[149]^x[129]^x[91]^x[80]^x[70]^x[64]^x[53]^x[47]^x[22]^x[21]^x[11]^x[10];
	y[20]=x[350]^x[341]^x[340]^x[330]^x[328]^x[314]^x[287]^x[276]^x[254]^x[248]^x[150]^x[148]^x[128]^x[94]^x[90]^x[84]^x[69]^x[52]^x[46]^x[30]^x[21]^x[20]^x[18]^x[10]^x[9];
	y[19]=x[349]^x[340]^x[339]^x[329]^x[327]^x[286]^x[275]^x[253]^x[247]^x[159]^x[149]^x[147]^x[138]^x[93]^x[51]^x[45]^x[29]^x[20]^x[19]^x[17]^x[9]^x[8];
	y[18]=x[348]^x[339]^x[338]^x[328]^x[326]^x[285]^x[274]^x[252]^x[246]^x[158]^x[148]^x[146]^x[137]^x[92]^x[50]^x[44]^x[28]^x[19]^x[18]^x[16]^x[8]^x[7];
	y[17]=x[347]^x[341]^x[338]^x[337]^x[335]^x[330]^x[327]^x[325]^x[324]^x[284]^x[273]^x[251]^x[245]^x[235]^x[234]^x[224]^x[181]^x[170]^x[157]^x[147]^x[145]^x[136]^x[91]^x[49]^x[43]^x[27]^x[18]^x[17]^x[15]^x[7]^x[6];
	y[16]=x[346]^x[340]^x[337]^x[336]^x[334]^x[329]^x[326]^x[324]^x[323]^x[283]^x[272]^x[250]^x[244]^x[233]^x[180]^x[169]^x[156]^x[146]^x[144]^x[135]^x[90]^x[48]^x[42]^x[26]^x[17]^x[16]^x[14]^x[6]^x[5];
	y[15]=x[345]^x[339]^x[336]^x[335]^x[333]^x[328]^x[325]^x[323]^x[322]^x[309]^x[298]^x[282]^x[271]^x[249]^x[243]^x[232]^x[179]^x[168]^x[155]^x[145]^x[143]^x[134]^x[89]^x[74]^x[68]^x[47]^x[41]^x[25]^x[16]^x[15]^x[13]^x[5]^x[4];
	y[14]=x[344]^x[338]^x[335]^x[334]^x[332]^x[327]^x[324]^x[322]^x[321]^x[308]^x[297]^x[281]^x[270]^x[248]^x[242]^x[231]^x[178]^x[167]^x[154]^x[144]^x[142]^x[133]^x[88]^x[73]^x[67]^x[46]^x[40]^x[24]^x[15]^x[14]^x[12]^x[4]^x[3];
	y[13]=x[343]^x[337]^x[334]^x[333]^x[331]^x[326]^x[323]^x[321]^x[320]^x[307]^x[296]^x[280]^x[269]^x[247]^x[241]^x[230]^x[177]^x[166]^x[153]^x[143]^x[141]^x[132]^x[87]^x[72]^x[66]^x[45]^x[39]^x[23]^x[14]^x[13]^x[11]^x[3]^x[2];
	y[12]=x[342]^x[336]^x[333]^x[332]^x[325]^x[322]^x[320]^x[306]^x[295]^x[279]^x[268]^x[246]^x[240]^x[229]^x[176]^x[165]^x[152]^x[142]^x[140]^x[131]^x[86]^x[71]^x[65]^x[44]^x[38]^x[22]^x[13]^x[12]^x[2]^x[1];
	y[11]=x[332]^x[331]^x[321]^x[305]^x[294]^x[278]^x[267]^x[235]^x[224]^x[151]^x[141]^x[139]^x[130]^x[75]^x[70]^x[43]^x[37]^x[12]^x[11]^x[1]^x[0];
	y[10]=x[331]^x[330]^x[320]^x[304]^x[293]^x[277]^x[266]^x[150]^x[140]^x[138]^x[129]^x[69]^x[42]^x[36]^x[11]^x[10]^x[0];
	y[9]=x[351]^x[329]^x[276]^x[265]^x[254]^x[248]^x[243]^x[237]^x[149]^x[139]^x[137]^x[128]^x[94]^x[83]^x[41]^x[35]^x[31]^x[19]^x[9]^x[7];
	y[8]=x[350]^x[328]^x[275]^x[264]^x[253]^x[247]^x[242]^x[236]^x[159]^x[148]^x[136]^x[93]^x[82]^x[40]^x[34]^x[30]^x[18]^x[8]^x[6];
	y[7]=x[349]^x[327]^x[274]^x[263]^x[252]^x[246]^x[241]^x[235]^x[158]^x[147]^x[135]^x[92]^x[81]^x[39]^x[33]^x[29]^x[17]^x[7]^x[5];
	y[6]=x[348]^x[326]^x[273]^x[262]^x[251]^x[245]^x[240]^x[234]^x[157]^x[146]^x[134]^x[91]^x[80]^x[38]^x[32]^x[28]^x[16]^x[6]^x[4];
	y[5]=x[347]^x[341]^x[335]^x[330]^x[325]^x[324]^x[310]^x[288]^x[272]^x[261]^x[250]^x[244]^x[239]^x[233]^x[181]^x[170]^x[156]^x[145]^x[133]^x[90]^x[79]^x[75]^x[69]^x[64]^x[37]^x[27]^x[15]^x[5]^x[3];
	y[4]=x[346]^x[340]^x[334]^x[329]^x[324]^x[323]^x[309]^x[298]^x[271]^x[260]^x[249]^x[243]^x[238]^x[232]^x[180]^x[169]^x[155]^x[144]^x[132]^x[89]^x[78]^x[74]^x[68]^x[36]^x[26]^x[14]^x[4]^x[2];
	y[3]=x[345]^x[339]^x[333]^x[328]^x[323]^x[322]^x[308]^x[297]^x[270]^x[259]^x[248]^x[242]^x[237]^x[231]^x[179]^x[168]^x[154]^x[143]^x[131]^x[88]^x[77]^x[73]^x[67]^x[35]^x[25]^x[13]^x[3]^x[1];
	y[2]=x[344]^x[338]^x[332]^x[327]^x[322]^x[321]^x[307]^x[296]^x[269]^x[258]^x[247]^x[241]^x[236]^x[230]^x[178]^x[167]^x[153]^x[142]^x[130]^x[87]^x[76]^x[72]^x[66]^x[34]^x[24]^x[12]^x[2]^x[0];
	y[1]=x[343]^x[337]^x[331]^x[326]^x[321]^x[320]^x[306]^x[295]^x[268]^x[257]^x[246]^x[240]^x[235]^x[229]^x[177]^x[166]^x[152]^x[141]^x[129]^x[86]^x[75]^x[71]^x[65]^x[33]^x[23]^x[11]^x[1];
	y[0]=x[342]^x[336]^x[325]^x[320]^x[305]^x[294]^x[267]^x[256]^x[176]^x[165]^x[151]^x[140]^x[128]^x[70]^x[64]^x[32]^x[22]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint44(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[381]^x[374]^x[372]^x[370]^x[363]^x[362]^x[359]^x[319]^x[317]^x[309]^x[308]^x[307]^x[299]^x[297]^x[295]^x[288]^x[282]^x[272]^x[261]^x[255]^x[245]^x[234]^x[223]^x[217]^x[212]^x[206]^x[159]^x[157]^x[153]^x[151]^x[149]^x[148]^x[143]^x[142]^x[139]^x[136]^x[135]^x[133]^x[130]^x[129]^x[128]^x[127]^x[108]^x[107]^x[97]^x[63]^x[58]^x[31]^x[25];
	y[30]=x[382]^x[380]^x[373]^x[370]^x[369]^x[362]^x[361]^x[359]^x[358]^x[319]^x[318]^x[316]^x[308]^x[307]^x[306]^x[296]^x[294]^x[254]^x[244]^x[233]^x[159]^x[158]^x[156]^x[153]^x[152]^x[150]^x[148]^x[142]^x[134]^x[128]^x[126]^x[107]^x[106]^x[96]^x[30]^x[24];
	y[29]=x[381]^x[379]^x[372]^x[369]^x[368]^x[361]^x[360]^x[358]^x[357]^x[318]^x[317]^x[315]^x[309]^x[307]^x[306]^x[305]^x[303]^x[298]^x[295]^x[293]^x[292]^x[253]^x[243]^x[232]^x[158]^x[157]^x[155]^x[152]^x[151]^x[147]^x[141]^x[138]^x[133]^x[127]^x[125]^x[105]^x[29]^x[23];
	y[28]=x[380]^x[378]^x[371]^x[368]^x[367]^x[360]^x[359]^x[357]^x[356]^x[317]^x[316]^x[314]^x[308]^x[306]^x[305]^x[304]^x[302]^x[297]^x[294]^x[292]^x[291]^x[252]^x[242]^x[231]^x[157]^x[156]^x[154]^x[151]^x[150]^x[146]^x[140]^x[137]^x[132]^x[126]^x[124]^x[104]^x[28]^x[22];
	y[27]=x[379]^x[377]^x[370]^x[367]^x[366]^x[359]^x[358]^x[356]^x[355]^x[316]^x[315]^x[313]^x[307]^x[305]^x[304]^x[303]^x[301]^x[296]^x[293]^x[291]^x[290]^x[251]^x[241]^x[230]^x[156]^x[155]^x[153]^x[150]^x[149]^x[145]^x[139]^x[136]^x[131]^x[125]^x[123]^x[103]^x[27]^x[21];
	y[26]=x[378]^x[376]^x[369]^x[366]^x[365]^x[358]^x[357]^x[355]^x[354]^x[319]^x[318]^x[315]^x[314]^x[313]^x[307]^x[304]^x[303]^x[302]^x[301]^x[292]^x[290]^x[277]^x[267]^x[256]^x[250]^x[240]^x[229]^x[212]^x[211]^x[201]^x[159]^x[158]^x[155]^x[154]^x[152]^x[149]^x[148]^x[147]^x[146]^x[144]^x[138]^x[130]^x[124]^x[122]^x[102]^x[53]^x[47]^x[26]^x[20];
	y[25]=x[377]^x[375]^x[368]^x[365]^x[364]^x[357]^x[356]^x[354]^x[353]^x[318]^x[317]^x[314]^x[313]^x[312]^x[306]^x[303]^x[302]^x[301]^x[300]^x[291]^x[289]^x[276]^x[249]^x[239]^x[228]^x[211]^x[210]^x[200]^x[158]^x[157]^x[154]^x[153]^x[151]^x[148]^x[147]^x[146]^x[145]^x[143]^x[137]^x[129]^x[123]^x[121]^x[101]^x[63]^x[57]^x[52]^x[46]^x[42]^x[36]^x[25]^x[19];
	y[24]=x[376]^x[374]^x[367]^x[364]^x[363]^x[356]^x[355]^x[353]^x[352]^x[317]^x[316]^x[313]^x[312]^x[311]^x[305]^x[302]^x[301]^x[300]^x[299]^x[290]^x[288]^x[275]^x[248]^x[238]^x[227]^x[210]^x[209]^x[199]^x[157]^x[156]^x[153]^x[152]^x[150]^x[147]^x[146]^x[145]^x[144]^x[142]^x[136]^x[128]^x[122]^x[120]^x[100]^x[62]^x[56]^x[51]^x[45]^x[41]^x[35]^x[24]^x[18];
	y[23]=x[375]^x[366]^x[355]^x[354]^x[316]^x[315]^x[312]^x[311]^x[310]^x[309]^x[304]^x[303]^x[301]^x[300]^x[299]^x[298]^x[292]^x[289]^x[274]^x[247]^x[237]^x[226]^x[209]^x[208]^x[198]^x[156]^x[155]^x[152]^x[151]^x[146]^x[145]^x[144]^x[143]^x[141]^x[135]^x[132]^x[121]^x[119]^x[99]^x[61]^x[55]^x[50]^x[44]^x[40]^x[34]^x[23]^x[17];
	y[22]=x[374]^x[365]^x[354]^x[353]^x[315]^x[314]^x[311]^x[310]^x[309]^x[308]^x[303]^x[302]^x[300]^x[299]^x[298]^x[297]^x[291]^x[288]^x[273]^x[246]^x[236]^x[225]^x[208]^x[207]^x[197]^x[155]^x[154]^x[151]^x[150]^x[145]^x[144]^x[143]^x[142]^x[140]^x[134]^x[131]^x[120]^x[118]^x[98]^x[60]^x[54]^x[49]^x[43]^x[39]^x[33]^x[22]^x[16];
	y[21]=x[364]^x[362]^x[353]^x[352]^x[314]^x[313]^x[310]^x[309]^x[308]^x[307]^x[302]^x[301]^x[299]^x[297]^x[296]^x[290]^x[272]^x[245]^x[235]^x[224]^x[213]^x[206]^x[202]^x[154]^x[153]^x[150]^x[149]^x[144]^x[143]^x[142]^x[141]^x[139]^x[138]^x[133]^x[132]^x[130]^x[119]^x[117]^x[97]^x[59]^x[48]^x[38]^x[32]^x[21]^x[15];
	y[20]=x[383]^x[382]^x[381]^x[372]^x[370]^x[363]^x[362]^x[352]^x[318]^x[309]^x[308]^x[298]^x[296]^x[282]^x[255]^x[244]^x[222]^x[216]^x[158]^x[152]^x[149]^x[148]^x[146]^x[143]^x[142]^x[140]^x[138]^x[137]^x[132]^x[131]^x[118]^x[116]^x[96]^x[62]^x[58]^x[52]^x[37]^x[20]^x[14];
	y[19]=x[383]^x[382]^x[381]^x[380]^x[371]^x[369]^x[361]^x[317]^x[308]^x[307]^x[297]^x[295]^x[254]^x[243]^x[221]^x[215]^x[157]^x[151]^x[148]^x[147]^x[145]^x[142]^x[141]^x[139]^x[137]^x[136]^x[131]^x[130]^x[127]^x[117]^x[115]^x[106]^x[61]^x[19]^x[13];
	y[18]=x[382]^x[381]^x[380]^x[379]^x[370]^x[368]^x[360]^x[316]^x[307]^x[306]^x[296]^x[294]^x[253]^x[242]^x[220]^x[214]^x[156]^x[150]^x[147]^x[146]^x[144]^x[141]^x[140]^x[138]^x[136]^x[135]^x[130]^x[129]^x[126]^x[116]^x[114]^x[105]^x[60]^x[18]^x[12];
	y[17]=x[381]^x[380]^x[379]^x[378]^x[369]^x[367]^x[359]^x[315]^x[309]^x[306]^x[305]^x[303]^x[298]^x[295]^x[293]^x[292]^x[252]^x[241]^x[219]^x[213]^x[203]^x[202]^x[192]^x[155]^x[146]^x[145]^x[143]^x[140]^x[139]^x[138]^x[137]^x[135]^x[134]^x[129]^x[128]^x[125]^x[115]^x[113]^x[104]^x[59]^x[17]^x[11];
	y[16]=x[380]^x[379]^x[378]^x[377]^x[368]^x[366]^x[358]^x[314]^x[308]^x[305]^x[304]^x[302]^x[297]^x[294]^x[292]^x[291]^x[251]^x[240]^x[218]^x[212]^x[201]^x[154]^x[145]^x[144]^x[142]^x[139]^x[138]^x[137]^x[136]^x[134]^x[133]^x[128]^x[124]^x[114]^x[112]^x[103]^x[58]^x[16]^x[10];
	y[15]=x[379]^x[378]^x[377]^x[376]^x[367]^x[365]^x[357]^x[313]^x[307]^x[304]^x[303]^x[301]^x[296]^x[293]^x[291]^x[290]^x[277]^x[266]^x[250]^x[239]^x[217]^x[211]^x[200]^x[153]^x[144]^x[143]^x[141]^x[138]^x[137]^x[136]^x[135]^x[133]^x[132]^x[123]^x[113]^x[111]^x[102]^x[57]^x[42]^x[36]^x[15]^x[9];
	y[14]=x[378]^x[377]^x[376]^x[375]^x[366]^x[364]^x[356]^x[312]^x[306]^x[303]^x[302]^x[300]^x[295]^x[292]^x[290]^x[289]^x[276]^x[265]^x[249]^x[238]^x[216]^x[210]^x[199]^x[152]^x[143]^x[142]^x[140]^x[137]^x[136]^x[135]^x[134]^x[132]^x[131]^x[122]^x[112]^x[110]^x[101]^x[56]^x[41]^x[35]^x[14]^x[8];
	y[13]=x[377]^x[376]^x[375]^x[374]^x[365]^x[363]^x[355]^x[311]^x[305]^x[302]^x[301]^x[299]^x[294]^x[291]^x[289]^x[288]^x[275]^x[264]^x[248]^x[237]^x[215]^x[209]^x[198]^x[151]^x[142]^x[141]^x[139]^x[136]^x[135]^x[134]^x[133]^x[131]^x[130]^x[121]^x[111]^x[109]^x[100]^x[55]^x[40]^x[34]^x[13]^x[7];
	y[12]=x[376]^x[375]^x[374]^x[364]^x[354]^x[310]^x[304]^x[301]^x[300]^x[293]^x[290]^x[288]^x[274]^x[263]^x[247]^x[236]^x[214]^x[208]^x[197]^x[150]^x[141]^x[140]^x[135]^x[134]^x[133]^x[130]^x[129]^x[120]^x[110]^x[108]^x[99]^x[54]^x[39]^x[33]^x[12]^x[6];
	y[11]=x[375]^x[374]^x[353]^x[352]^x[300]^x[299]^x[289]^x[273]^x[262]^x[246]^x[235]^x[203]^x[192]^x[140]^x[139]^x[134]^x[133]^x[129]^x[128]^x[119]^x[109]^x[107]^x[98]^x[43]^x[38]^x[11]^x[5];
	y[10]=x[374]^x[373]^x[362]^x[352]^x[299]^x[298]^x[288]^x[272]^x[261]^x[245]^x[234]^x[139]^x[138]^x[133]^x[132]^x[128]^x[118]^x[108]^x[106]^x[97]^x[37]^x[10]^x[4];
	y[9]=x[383]^x[382]^x[373]^x[372]^x[371]^x[370]^x[362]^x[361]^x[359]^x[319]^x[297]^x[244]^x[233]^x[222]^x[216]^x[211]^x[205]^x[159]^x[153]^x[147]^x[141]^x[137]^x[135]^x[131]^x[129]^x[117]^x[107]^x[105]^x[96]^x[62]^x[51]^x[9]^x[3];
	y[8]=x[382]^x[381]^x[372]^x[371]^x[370]^x[369]^x[361]^x[360]^x[358]^x[318]^x[296]^x[243]^x[232]^x[221]^x[215]^x[210]^x[204]^x[158]^x[152]^x[146]^x[140]^x[136]^x[134]^x[130]^x[128]^x[127]^x[116]^x[104]^x[61]^x[50]^x[8]^x[2];
	y[7]=x[381]^x[380]^x[371]^x[370]^x[369]^x[368]^x[360]^x[359]^x[357]^x[317]^x[295]^x[242]^x[231]^x[220]^x[214]^x[209]^x[203]^x[157]^x[151]^x[145]^x[139]^x[135]^x[133]^x[129]^x[126]^x[115]^x[103]^x[60]^x[49]^x[7]^x[1];
	y[6]=x[380]^x[379]^x[370]^x[369]^x[368]^x[367]^x[359]^x[358]^x[356]^x[316]^x[294]^x[241]^x[230]^x[219]^x[213]^x[208]^x[202]^x[156]^x[150]^x[144]^x[138]^x[134]^x[132]^x[128]^x[125]^x[114]^x[102]^x[59]^x[48]^x[6]^x[0];
	y[5]=x[379]^x[378]^x[369]^x[368]^x[367]^x[366]^x[358]^x[357]^x[355]^x[315]^x[309]^x[303]^x[298]^x[293]^x[292]^x[278]^x[256]^x[240]^x[229]^x[218]^x[212]^x[207]^x[201]^x[155]^x[143]^x[138]^x[137]^x[133]^x[131]^x[124]^x[113]^x[101]^x[58]^x[47]^x[43]^x[37]^x[32]^x[5];
	y[4]=x[378]^x[377]^x[368]^x[367]^x[366]^x[365]^x[357]^x[356]^x[354]^x[314]^x[308]^x[302]^x[297]^x[292]^x[291]^x[277]^x[266]^x[239]^x[228]^x[217]^x[211]^x[206]^x[200]^x[154]^x[142]^x[137]^x[136]^x[132]^x[130]^x[123]^x[112]^x[100]^x[57]^x[46]^x[42]^x[36]^x[4];
	y[3]=x[377]^x[376]^x[367]^x[366]^x[365]^x[364]^x[356]^x[355]^x[353]^x[313]^x[307]^x[301]^x[296]^x[291]^x[290]^x[276]^x[265]^x[238]^x[227]^x[216]^x[210]^x[205]^x[199]^x[153]^x[141]^x[136]^x[135]^x[131]^x[129]^x[122]^x[111]^x[99]^x[56]^x[45]^x[41]^x[35]^x[3];
	y[2]=x[376]^x[375]^x[366]^x[365]^x[364]^x[363]^x[355]^x[354]^x[352]^x[312]^x[306]^x[300]^x[295]^x[290]^x[289]^x[275]^x[264]^x[237]^x[226]^x[215]^x[209]^x[204]^x[198]^x[152]^x[140]^x[135]^x[134]^x[130]^x[128]^x[121]^x[110]^x[98]^x[55]^x[44]^x[40]^x[34]^x[2];
	y[1]=x[375]^x[374]^x[365]^x[364]^x[363]^x[354]^x[353]^x[311]^x[305]^x[299]^x[294]^x[289]^x[288]^x[274]^x[263]^x[236]^x[225]^x[214]^x[208]^x[203]^x[197]^x[151]^x[139]^x[134]^x[133]^x[129]^x[120]^x[109]^x[97]^x[54]^x[43]^x[39]^x[33]^x[1];
	y[0]=x[374]^x[364]^x[363]^x[353]^x[352]^x[310]^x[304]^x[293]^x[288]^x[273]^x[262]^x[235]^x[224]^x[150]^x[133]^x[128]^x[119]^x[108]^x[96]^x[38]^x[32]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint45(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[377]^x[373]^x[367]^x[362]^x[356]^x[349]^x[342]^x[340]^x[338]^x[331]^x[330]^x[327]^x[287]^x[285]^x[277]^x[276]^x[275]^x[267]^x[265]^x[263]^x[256]^x[250]^x[240]^x[229]^x[223]^x[213]^x[202]^x[191]^x[185]^x[180]^x[174]^x[159]^x[147]^x[127]^x[125]^x[121]^x[119]^x[117]^x[116]^x[111]^x[110]^x[107]^x[104]^x[103]^x[101]^x[98]^x[97]^x[96]^x[95]^x[76]^x[75]^x[65]^x[31]^x[26];
	y[30]=x[382]^x[376]^x[372]^x[366]^x[361]^x[355]^x[350]^x[348]^x[341]^x[338]^x[337]^x[330]^x[329]^x[327]^x[326]^x[287]^x[286]^x[284]^x[276]^x[275]^x[274]^x[264]^x[262]^x[222]^x[212]^x[201]^x[158]^x[146]^x[127]^x[126]^x[124]^x[121]^x[120]^x[118]^x[116]^x[110]^x[102]^x[96]^x[94]^x[75]^x[74]^x[64];
	y[29]=x[381]^x[375]^x[371]^x[365]^x[360]^x[354]^x[349]^x[347]^x[340]^x[337]^x[336]^x[329]^x[328]^x[326]^x[325]^x[286]^x[285]^x[283]^x[277]^x[275]^x[274]^x[273]^x[271]^x[266]^x[263]^x[261]^x[260]^x[221]^x[211]^x[200]^x[157]^x[145]^x[126]^x[125]^x[123]^x[120]^x[119]^x[115]^x[109]^x[106]^x[101]^x[95]^x[93]^x[73];
	y[28]=x[380]^x[374]^x[370]^x[364]^x[359]^x[353]^x[348]^x[346]^x[339]^x[336]^x[335]^x[328]^x[327]^x[325]^x[324]^x[285]^x[284]^x[282]^x[276]^x[274]^x[273]^x[272]^x[270]^x[265]^x[262]^x[260]^x[259]^x[220]^x[210]^x[199]^x[156]^x[144]^x[125]^x[124]^x[122]^x[119]^x[118]^x[114]^x[108]^x[105]^x[100]^x[94]^x[92]^x[72];
	y[27]=x[379]^x[373]^x[369]^x[363]^x[358]^x[352]^x[347]^x[345]^x[338]^x[335]^x[334]^x[327]^x[326]^x[324]^x[323]^x[284]^x[283]^x[281]^x[275]^x[273]^x[272]^x[271]^x[269]^x[264]^x[261]^x[259]^x[258]^x[219]^x[209]^x[198]^x[155]^x[143]^x[124]^x[123]^x[121]^x[118]^x[117]^x[113]^x[107]^x[104]^x[99]^x[93]^x[91]^x[71];
	y[26]=x[383]^x[378]^x[372]^x[368]^x[357]^x[346]^x[344]^x[337]^x[334]^x[333]^x[326]^x[325]^x[323]^x[322]^x[287]^x[286]^x[283]^x[282]^x[281]^x[275]^x[272]^x[271]^x[270]^x[269]^x[260]^x[258]^x[245]^x[235]^x[224]^x[218]^x[208]^x[197]^x[180]^x[179]^x[169]^x[154]^x[142]^x[127]^x[126]^x[123]^x[122]^x[120]^x[117]^x[116]^x[115]^x[114]^x[112]^x[106]^x[98]^x[92]^x[90]^x[70]^x[21]^x[15];
	y[25]=x[382]^x[377]^x[371]^x[367]^x[356]^x[345]^x[343]^x[336]^x[333]^x[332]^x[325]^x[324]^x[322]^x[321]^x[286]^x[285]^x[282]^x[281]^x[280]^x[274]^x[271]^x[270]^x[269]^x[268]^x[259]^x[257]^x[244]^x[217]^x[207]^x[196]^x[179]^x[178]^x[168]^x[153]^x[141]^x[126]^x[125]^x[122]^x[121]^x[119]^x[116]^x[115]^x[114]^x[113]^x[111]^x[105]^x[97]^x[91]^x[89]^x[69]^x[31]^x[25]^x[20]^x[14]^x[10]^x[4];
	y[24]=x[381]^x[376]^x[370]^x[366]^x[355]^x[344]^x[342]^x[335]^x[332]^x[331]^x[324]^x[323]^x[321]^x[320]^x[285]^x[284]^x[281]^x[280]^x[279]^x[273]^x[270]^x[269]^x[268]^x[267]^x[258]^x[256]^x[243]^x[216]^x[206]^x[195]^x[178]^x[177]^x[167]^x[152]^x[140]^x[125]^x[124]^x[121]^x[120]^x[118]^x[115]^x[114]^x[113]^x[112]^x[110]^x[104]^x[96]^x[90]^x[88]^x[68]^x[30]^x[24]^x[19]^x[13]^x[9]^x[3];
	y[23]=x[380]^x[375]^x[369]^x[365]^x[354]^x[343]^x[334]^x[323]^x[322]^x[284]^x[283]^x[280]^x[279]^x[278]^x[277]^x[272]^x[271]^x[269]^x[268]^x[267]^x[266]^x[260]^x[257]^x[242]^x[215]^x[205]^x[194]^x[177]^x[176]^x[166]^x[151]^x[139]^x[124]^x[123]^x[120]^x[119]^x[114]^x[113]^x[112]^x[111]^x[109]^x[103]^x[100]^x[89]^x[87]^x[67]^x[29]^x[23]^x[18]^x[12]^x[8]^x[2];
	y[22]=x[379]^x[374]^x[368]^x[364]^x[353]^x[342]^x[333]^x[322]^x[321]^x[283]^x[282]^x[279]^x[278]^x[277]^x[276]^x[271]^x[270]^x[268]^x[267]^x[266]^x[265]^x[259]^x[256]^x[241]^x[214]^x[204]^x[193]^x[176]^x[175]^x[165]^x[150]^x[138]^x[123]^x[122]^x[119]^x[118]^x[113]^x[112]^x[111]^x[110]^x[108]^x[102]^x[99]^x[88]^x[86]^x[66]^x[28]^x[22]^x[17]^x[11]^x[7]^x[1];
	y[21]=x[378]^x[373]^x[367]^x[363]^x[352]^x[332]^x[330]^x[321]^x[320]^x[282]^x[281]^x[278]^x[277]^x[276]^x[275]^x[270]^x[269]^x[267]^x[265]^x[264]^x[258]^x[240]^x[213]^x[203]^x[192]^x[181]^x[174]^x[170]^x[149]^x[137]^x[122]^x[121]^x[118]^x[117]^x[112]^x[111]^x[110]^x[109]^x[107]^x[106]^x[101]^x[100]^x[98]^x[87]^x[85]^x[65]^x[27]^x[16]^x[6]^x[0];
	y[20]=x[383]^x[377]^x[372]^x[366]^x[351]^x[350]^x[349]^x[340]^x[338]^x[331]^x[330]^x[320]^x[286]^x[277]^x[276]^x[266]^x[264]^x[250]^x[223]^x[212]^x[190]^x[184]^x[148]^x[136]^x[126]^x[120]^x[117]^x[116]^x[114]^x[111]^x[110]^x[108]^x[106]^x[105]^x[100]^x[99]^x[86]^x[84]^x[64]^x[30]^x[26]^x[20]^x[5];
	y[19]=x[382]^x[376]^x[371]^x[365]^x[351]^x[350]^x[349]^x[348]^x[339]^x[337]^x[329]^x[285]^x[276]^x[275]^x[265]^x[263]^x[222]^x[211]^x[189]^x[183]^x[147]^x[135]^x[125]^x[119]^x[116]^x[115]^x[113]^x[110]^x[109]^x[107]^x[105]^x[104]^x[99]^x[98]^x[95]^x[85]^x[83]^x[74]^x[29];
	y[18]=x[381]^x[375]^x[370]^x[364]^x[350]^x[349]^x[348]^x[347]^x[338]^x[336]^x[328]^x[284]^x[275]^x[274]^x[264]^x[262]^x[221]^x[210]^x[188]^x[182]^x[146]^x[134]^x[124]^x[118]^x[115]^x[114]^x[112]^x[109]^x[108]^x[106]^x[104]^x[103]^x[98]^x[97]^x[94]^x[84]^x[82]^x[73]^x[28];
	y[17]=x[380]^x[374]^x[369]^x[363]^x[349]^x[348]^x[347]^x[346]^x[337]^x[335]^x[327]^x[283]^x[277]^x[274]^x[273]^x[271]^x[266]^x[263]^x[261]^x[260]^x[220]^x[209]^x[187]^x[181]^x[171]^x[170]^x[160]^x[145]^x[133]^x[123]^x[114]^x[113]^x[111]^x[108]^x[107]^x[106]^x[105]^x[103]^x[102]^x[97]^x[96]^x[93]^x[83]^x[81]^x[72]^x[27];
	y[16]=x[379]^x[373]^x[368]^x[362]^x[348]^x[347]^x[346]^x[345]^x[336]^x[334]^x[326]^x[282]^x[276]^x[273]^x[272]^x[270]^x[265]^x[262]^x[260]^x[259]^x[219]^x[208]^x[186]^x[180]^x[169]^x[144]^x[132]^x[122]^x[113]^x[112]^x[110]^x[107]^x[106]^x[105]^x[104]^x[102]^x[101]^x[96]^x[92]^x[82]^x[80]^x[71]^x[26];
	y[15]=x[378]^x[372]^x[367]^x[361]^x[347]^x[346]^x[345]^x[344]^x[335]^x[333]^x[325]^x[281]^x[275]^x[272]^x[271]^x[269]^x[264]^x[261]^x[259]^x[258]^x[245]^x[234]^x[218]^x[207]^x[185]^x[179]^x[168]^x[143]^x[131]^x[121]^x[112]^x[111]^x[109]^x[106]^x[105]^x[104]^x[103]^x[101]^x[100]^x[91]^x[81]^x[79]^x[70]^x[25]^x[10]^x[4];
	y[14]=x[377]^x[371]^x[366]^x[360]^x[346]^x[345]^x[344]^x[343]^x[334]^x[332]^x[324]^x[280]^x[274]^x[271]^x[270]^x[268]^x[263]^x[260]^x[258]^x[257]^x[244]^x[233]^x[217]^x[206]^x[184]^x[178]^x[167]^x[142]^x[130]^x[120]^x[111]^x[110]^x[108]^x[105]^x[104]^x[103]^x[102]^x[100]^x[99]^x[90]^x[80]^x[78]^x[69]^x[24]^x[9]^x[3];
	y[13]=x[376]^x[370]^x[365]^x[359]^x[345]^x[344]^x[343]^x[342]^x[333]^x[331]^x[323]^x[279]^x[273]^x[270]^x[269]^x[267]^x[262]^x[259]^x[257]^x[256]^x[243]^x[232]^x[216]^x[205]^x[183]^x[177]^x[166]^x[141]^x[129]^x[119]^x[110]^x[109]^x[107]^x[104]^x[103]^x[102]^x[101]^x[99]^x[98]^x[89]^x[79]^x[77]^x[68]^x[23]^x[8]^x[2];
	y[12]=x[375]^x[369]^x[364]^x[358]^x[344]^x[343]^x[342]^x[332]^x[322]^x[278]^x[272]^x[269]^x[268]^x[261]^x[258]^x[256]^x[242]^x[231]^x[215]^x[204]^x[182]^x[176]^x[165]^x[140]^x[128]^x[118]^x[109]^x[108]^x[103]^x[102]^x[101]^x[98]^x[97]^x[88]^x[78]^x[76]^x[67]^x[22]^x[7]^x[1];
	y[11]=x[374]^x[368]^x[363]^x[357]^x[343]^x[342]^x[321]^x[320]^x[268]^x[267]^x[257]^x[241]^x[230]^x[214]^x[203]^x[171]^x[160]^x[139]^x[108]^x[107]^x[102]^x[101]^x[97]^x[96]^x[87]^x[77]^x[75]^x[66]^x[11]^x[6];
	y[10]=x[373]^x[367]^x[362]^x[356]^x[342]^x[341]^x[330]^x[320]^x[267]^x[266]^x[256]^x[240]^x[229]^x[213]^x[202]^x[138]^x[107]^x[106]^x[101]^x[100]^x[96]^x[86]^x[76]^x[74]^x[65]^x[5];
	y[9]=x[372]^x[366]^x[361]^x[355]^x[351]^x[350]^x[341]^x[340]^x[339]^x[338]^x[330]^x[329]^x[327]^x[287]^x[265]^x[212]^x[201]^x[190]^x[184]^x[179]^x[173]^x[137]^x[127]^x[121]^x[115]^x[109]^x[105]^x[103]^x[99]^x[97]^x[85]^x[75]^x[73]^x[64]^x[30]^x[19];
	y[8]=x[371]^x[365]^x[360]^x[354]^x[350]^x[349]^x[340]^x[339]^x[338]^x[337]^x[329]^x[328]^x[326]^x[286]^x[264]^x[211]^x[200]^x[189]^x[183]^x[178]^x[172]^x[136]^x[126]^x[120]^x[114]^x[108]^x[104]^x[102]^x[98]^x[96]^x[95]^x[84]^x[72]^x[29]^x[18];
	y[7]=x[370]^x[364]^x[359]^x[353]^x[349]^x[348]^x[339]^x[338]^x[337]^x[336]^x[328]^x[327]^x[325]^x[285]^x[263]^x[210]^x[199]^x[188]^x[182]^x[177]^x[171]^x[135]^x[125]^x[119]^x[113]^x[107]^x[103]^x[101]^x[97]^x[94]^x[83]^x[71]^x[28]^x[17];
	y[6]=x[369]^x[363]^x[358]^x[352]^x[348]^x[347]^x[338]^x[337]^x[336]^x[335]^x[327]^x[326]^x[324]^x[284]^x[262]^x[209]^x[198]^x[187]^x[181]^x[176]^x[170]^x[134]^x[124]^x[118]^x[112]^x[106]^x[102]^x[100]^x[96]^x[93]^x[82]^x[70]^x[27]^x[16];
	y[5]=x[368]^x[357]^x[347]^x[346]^x[337]^x[336]^x[335]^x[334]^x[326]^x[325]^x[323]^x[283]^x[277]^x[271]^x[266]^x[261]^x[260]^x[246]^x[224]^x[208]^x[197]^x[186]^x[180]^x[175]^x[169]^x[133]^x[123]^x[111]^x[106]^x[105]^x[101]^x[99]^x[92]^x[81]^x[69]^x[26]^x[15]^x[11]^x[5]^x[0];
	y[4]=x[367]^x[356]^x[346]^x[345]^x[336]^x[335]^x[334]^x[333]^x[325]^x[324]^x[322]^x[282]^x[276]^x[270]^x[265]^x[260]^x[259]^x[245]^x[234]^x[207]^x[196]^x[185]^x[179]^x[174]^x[168]^x[132]^x[122]^x[110]^x[105]^x[104]^x[100]^x[98]^x[91]^x[80]^x[68]^x[25]^x[14]^x[10]^x[4];
	y[3]=x[366]^x[355]^x[345]^x[344]^x[335]^x[334]^x[333]^x[332]^x[324]^x[323]^x[321]^x[281]^x[275]^x[269]^x[264]^x[259]^x[258]^x[244]^x[233]^x[206]^x[195]^x[184]^x[178]^x[173]^x[167]^x[131]^x[121]^x[109]^x[104]^x[103]^x[99]^x[97]^x[90]^x[79]^x[67]^x[24]^x[13]^x[9]^x[3];
	y[2]=x[365]^x[354]^x[344]^x[343]^x[334]^x[333]^x[332]^x[331]^x[323]^x[322]^x[320]^x[280]^x[274]^x[268]^x[263]^x[258]^x[257]^x[243]^x[232]^x[205]^x[194]^x[183]^x[177]^x[172]^x[166]^x[130]^x[120]^x[108]^x[103]^x[102]^x[98]^x[96]^x[89]^x[78]^x[66]^x[23]^x[12]^x[8]^x[2];
	y[1]=x[364]^x[353]^x[343]^x[342]^x[333]^x[332]^x[331]^x[322]^x[321]^x[279]^x[273]^x[267]^x[262]^x[257]^x[256]^x[242]^x[231]^x[204]^x[193]^x[182]^x[176]^x[171]^x[165]^x[129]^x[119]^x[107]^x[102]^x[101]^x[97]^x[88]^x[77]^x[65]^x[22]^x[11]^x[7]^x[1];
	y[0]=x[363]^x[352]^x[342]^x[332]^x[331]^x[321]^x[320]^x[278]^x[272]^x[261]^x[256]^x[241]^x[230]^x[203]^x[192]^x[128]^x[118]^x[101]^x[96]^x[87]^x[76]^x[64]^x[6]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint46(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[378]^x[373]^x[368]^x[362]^x[357]^x[351]^x[345]^x[341]^x[335]^x[330]^x[324]^x[317]^x[310]^x[308]^x[306]^x[299]^x[298]^x[295]^x[255]^x[253]^x[245]^x[244]^x[243]^x[235]^x[233]^x[231]^x[224]^x[218]^x[208]^x[197]^x[191]^x[181]^x[170]^x[154]^x[142]^x[127]^x[115]^x[95]^x[93]^x[89]^x[87]^x[85]^x[84]^x[79]^x[78]^x[75]^x[72]^x[71]^x[69]^x[66]^x[65]^x[64]^x[63]^x[44]^x[43]^x[33];
	y[30]=x[350]^x[344]^x[340]^x[334]^x[329]^x[323]^x[318]^x[316]^x[309]^x[306]^x[305]^x[298]^x[297]^x[295]^x[294]^x[255]^x[254]^x[252]^x[244]^x[243]^x[242]^x[232]^x[230]^x[190]^x[180]^x[169]^x[126]^x[114]^x[95]^x[94]^x[92]^x[89]^x[88]^x[86]^x[84]^x[78]^x[70]^x[64]^x[62]^x[43]^x[42]^x[32];
	y[29]=x[349]^x[343]^x[339]^x[333]^x[328]^x[322]^x[317]^x[315]^x[308]^x[305]^x[304]^x[297]^x[296]^x[294]^x[293]^x[254]^x[253]^x[251]^x[245]^x[243]^x[242]^x[241]^x[239]^x[234]^x[231]^x[229]^x[228]^x[189]^x[179]^x[168]^x[125]^x[113]^x[94]^x[93]^x[91]^x[88]^x[87]^x[83]^x[77]^x[74]^x[69]^x[63]^x[61]^x[41];
	y[28]=x[348]^x[342]^x[338]^x[332]^x[327]^x[321]^x[316]^x[314]^x[307]^x[304]^x[303]^x[296]^x[295]^x[293]^x[292]^x[253]^x[252]^x[250]^x[244]^x[242]^x[241]^x[240]^x[238]^x[233]^x[230]^x[228]^x[227]^x[188]^x[178]^x[167]^x[124]^x[112]^x[93]^x[92]^x[90]^x[87]^x[86]^x[82]^x[76]^x[73]^x[68]^x[62]^x[60]^x[40];
	y[27]=x[347]^x[341]^x[337]^x[331]^x[326]^x[320]^x[315]^x[313]^x[306]^x[303]^x[302]^x[295]^x[294]^x[292]^x[291]^x[252]^x[251]^x[249]^x[243]^x[241]^x[240]^x[239]^x[237]^x[232]^x[229]^x[227]^x[226]^x[187]^x[177]^x[166]^x[123]^x[111]^x[92]^x[91]^x[89]^x[86]^x[85]^x[81]^x[75]^x[72]^x[67]^x[61]^x[59]^x[39];
	y[26]=x[378]^x[373]^x[367]^x[363]^x[352]^x[351]^x[346]^x[340]^x[336]^x[325]^x[314]^x[312]^x[305]^x[302]^x[301]^x[294]^x[293]^x[291]^x[290]^x[255]^x[254]^x[251]^x[250]^x[249]^x[243]^x[240]^x[239]^x[238]^x[237]^x[228]^x[226]^x[213]^x[203]^x[192]^x[186]^x[176]^x[165]^x[149]^x[148]^x[147]^x[122]^x[110]^x[95]^x[94]^x[91]^x[90]^x[88]^x[85]^x[84]^x[83]^x[82]^x[80]^x[74]^x[66]^x[60]^x[58]^x[38];
	y[25]=x[372]^x[366]^x[350]^x[345]^x[339]^x[335]^x[324]^x[313]^x[311]^x[304]^x[301]^x[300]^x[293]^x[292]^x[290]^x[289]^x[254]^x[253]^x[250]^x[249]^x[248]^x[242]^x[239]^x[238]^x[237]^x[236]^x[227]^x[225]^x[212]^x[185]^x[175]^x[164]^x[159]^x[148]^x[146]^x[138]^x[121]^x[109]^x[94]^x[93]^x[90]^x[89]^x[87]^x[84]^x[83]^x[82]^x[81]^x[79]^x[73]^x[65]^x[59]^x[57]^x[37];
	y[24]=x[371]^x[365]^x[349]^x[344]^x[338]^x[334]^x[323]^x[312]^x[310]^x[303]^x[300]^x[299]^x[292]^x[291]^x[289]^x[288]^x[253]^x[252]^x[249]^x[248]^x[247]^x[241]^x[238]^x[237]^x[236]^x[235]^x[226]^x[224]^x[211]^x[184]^x[174]^x[163]^x[158]^x[147]^x[145]^x[137]^x[120]^x[108]^x[93]^x[92]^x[89]^x[88]^x[86]^x[83]^x[82]^x[81]^x[80]^x[78]^x[72]^x[64]^x[58]^x[56]^x[36];
	y[23]=x[370]^x[364]^x[348]^x[343]^x[337]^x[333]^x[322]^x[311]^x[302]^x[291]^x[290]^x[252]^x[251]^x[248]^x[247]^x[246]^x[245]^x[240]^x[239]^x[237]^x[236]^x[235]^x[234]^x[228]^x[225]^x[210]^x[183]^x[173]^x[162]^x[157]^x[146]^x[144]^x[136]^x[119]^x[107]^x[92]^x[91]^x[88]^x[87]^x[82]^x[81]^x[80]^x[79]^x[77]^x[71]^x[68]^x[57]^x[55]^x[35];
	y[22]=x[369]^x[363]^x[347]^x[342]^x[336]^x[332]^x[321]^x[310]^x[301]^x[290]^x[289]^x[251]^x[250]^x[247]^x[246]^x[245]^x[244]^x[239]^x[238]^x[236]^x[235]^x[234]^x[233]^x[227]^x[224]^x[209]^x[182]^x[172]^x[161]^x[156]^x[145]^x[143]^x[135]^x[118]^x[106]^x[91]^x[90]^x[87]^x[86]^x[81]^x[80]^x[79]^x[78]^x[76]^x[70]^x[67]^x[56]^x[54]^x[34];
	y[21]=x[368]^x[363]^x[352]^x[346]^x[341]^x[335]^x[331]^x[320]^x[300]^x[298]^x[289]^x[288]^x[250]^x[249]^x[246]^x[245]^x[244]^x[243]^x[238]^x[237]^x[235]^x[233]^x[232]^x[226]^x[208]^x[181]^x[171]^x[160]^x[155]^x[144]^x[142]^x[134]^x[117]^x[105]^x[90]^x[89]^x[86]^x[85]^x[80]^x[79]^x[78]^x[77]^x[75]^x[74]^x[69]^x[68]^x[66]^x[55]^x[53]^x[33];
	y[20]=x[383]^x[382]^x[378]^x[361]^x[351]^x[345]^x[340]^x[334]^x[319]^x[318]^x[317]^x[308]^x[306]^x[299]^x[298]^x[288]^x[254]^x[245]^x[244]^x[234]^x[232]^x[218]^x[191]^x[180]^x[154]^x[142]^x[133]^x[116]^x[104]^x[94]^x[88]^x[85]^x[84]^x[82]^x[79]^x[78]^x[76]^x[74]^x[73]^x[68]^x[67]^x[54]^x[52]^x[32];
	y[19]=x[381]^x[371]^x[360]^x[350]^x[344]^x[339]^x[333]^x[319]^x[318]^x[317]^x[316]^x[307]^x[305]^x[297]^x[253]^x[244]^x[243]^x[233]^x[231]^x[190]^x[179]^x[115]^x[103]^x[93]^x[87]^x[84]^x[83]^x[81]^x[78]^x[77]^x[75]^x[73]^x[72]^x[67]^x[66]^x[63]^x[53]^x[51]^x[42];
	y[18]=x[380]^x[370]^x[359]^x[349]^x[343]^x[338]^x[332]^x[318]^x[317]^x[316]^x[315]^x[306]^x[304]^x[296]^x[252]^x[243]^x[242]^x[232]^x[230]^x[189]^x[178]^x[114]^x[102]^x[92]^x[86]^x[83]^x[82]^x[80]^x[77]^x[76]^x[74]^x[72]^x[71]^x[66]^x[65]^x[62]^x[52]^x[50]^x[41];
	y[17]=x[379]^x[369]^x[358]^x[348]^x[342]^x[337]^x[331]^x[317]^x[316]^x[315]^x[314]^x[305]^x[303]^x[295]^x[251]^x[245]^x[242]^x[241]^x[239]^x[234]^x[231]^x[229]^x[228]^x[188]^x[177]^x[139]^x[138]^x[128]^x[113]^x[101]^x[91]^x[82]^x[81]^x[79]^x[76]^x[75]^x[74]^x[73]^x[71]^x[70]^x[65]^x[64]^x[61]^x[51]^x[49]^x[40];
	y[16]=x[378]^x[368]^x[357]^x[347]^x[341]^x[336]^x[330]^x[316]^x[315]^x[314]^x[313]^x[304]^x[302]^x[294]^x[250]^x[244]^x[241]^x[240]^x[238]^x[233]^x[230]^x[228]^x[227]^x[187]^x[176]^x[137]^x[112]^x[100]^x[90]^x[81]^x[80]^x[78]^x[75]^x[74]^x[73]^x[72]^x[70]^x[69]^x[64]^x[60]^x[50]^x[48]^x[39];
	y[15]=x[377]^x[373]^x[362]^x[346]^x[340]^x[335]^x[329]^x[315]^x[314]^x[313]^x[312]^x[303]^x[301]^x[293]^x[249]^x[243]^x[240]^x[239]^x[237]^x[232]^x[229]^x[227]^x[226]^x[213]^x[202]^x[186]^x[175]^x[138]^x[136]^x[111]^x[99]^x[89]^x[80]^x[79]^x[77]^x[74]^x[73]^x[72]^x[71]^x[69]^x[68]^x[59]^x[49]^x[47]^x[38];
	y[14]=x[376]^x[372]^x[361]^x[345]^x[339]^x[334]^x[328]^x[314]^x[313]^x[312]^x[311]^x[302]^x[300]^x[292]^x[248]^x[242]^x[239]^x[238]^x[236]^x[231]^x[228]^x[226]^x[225]^x[212]^x[201]^x[185]^x[174]^x[137]^x[135]^x[110]^x[98]^x[88]^x[79]^x[78]^x[76]^x[73]^x[72]^x[71]^x[70]^x[68]^x[67]^x[58]^x[48]^x[46]^x[37];
	y[13]=x[375]^x[371]^x[360]^x[344]^x[338]^x[333]^x[327]^x[313]^x[312]^x[311]^x[310]^x[301]^x[299]^x[291]^x[247]^x[241]^x[238]^x[237]^x[235]^x[230]^x[227]^x[225]^x[224]^x[211]^x[200]^x[184]^x[173]^x[136]^x[134]^x[109]^x[97]^x[87]^x[78]^x[77]^x[75]^x[72]^x[71]^x[70]^x[69]^x[67]^x[66]^x[57]^x[47]^x[45]^x[36];
	y[12]=x[374]^x[370]^x[359]^x[343]^x[337]^x[332]^x[326]^x[312]^x[311]^x[310]^x[300]^x[290]^x[246]^x[240]^x[237]^x[236]^x[229]^x[226]^x[224]^x[210]^x[199]^x[183]^x[172]^x[135]^x[133]^x[108]^x[96]^x[86]^x[77]^x[76]^x[71]^x[70]^x[69]^x[66]^x[65]^x[56]^x[46]^x[44]^x[35];
	y[11]=x[374]^x[369]^x[363]^x[358]^x[342]^x[336]^x[331]^x[325]^x[311]^x[310]^x[289]^x[288]^x[236]^x[235]^x[225]^x[209]^x[198]^x[182]^x[171]^x[134]^x[133]^x[107]^x[76]^x[75]^x[70]^x[69]^x[65]^x[64]^x[55]^x[45]^x[43]^x[34];
	y[10]=x[368]^x[357]^x[341]^x[335]^x[330]^x[324]^x[310]^x[309]^x[298]^x[288]^x[235]^x[234]^x[224]^x[208]^x[197]^x[181]^x[170]^x[133]^x[106]^x[75]^x[74]^x[69]^x[68]^x[64]^x[54]^x[44]^x[42]^x[33];
	y[9]=x[372]^x[371]^x[361]^x[340]^x[334]^x[329]^x[323]^x[319]^x[318]^x[309]^x[308]^x[307]^x[306]^x[298]^x[297]^x[295]^x[255]^x[233]^x[180]^x[169]^x[105]^x[95]^x[89]^x[83]^x[77]^x[73]^x[71]^x[67]^x[65]^x[53]^x[43]^x[41]^x[32];
	y[8]=x[371]^x[370]^x[360]^x[339]^x[333]^x[328]^x[322]^x[318]^x[317]^x[308]^x[307]^x[306]^x[305]^x[297]^x[296]^x[294]^x[254]^x[232]^x[179]^x[168]^x[104]^x[94]^x[88]^x[82]^x[76]^x[72]^x[70]^x[66]^x[64]^x[63]^x[52]^x[40];
	y[7]=x[370]^x[369]^x[359]^x[338]^x[332]^x[327]^x[321]^x[317]^x[316]^x[307]^x[306]^x[305]^x[304]^x[296]^x[295]^x[293]^x[253]^x[231]^x[178]^x[167]^x[103]^x[93]^x[87]^x[81]^x[75]^x[71]^x[69]^x[65]^x[62]^x[51]^x[39];
	y[6]=x[369]^x[368]^x[358]^x[337]^x[331]^x[326]^x[320]^x[316]^x[315]^x[306]^x[305]^x[304]^x[303]^x[295]^x[294]^x[292]^x[252]^x[230]^x[177]^x[166]^x[102]^x[92]^x[86]^x[80]^x[74]^x[70]^x[68]^x[64]^x[61]^x[50]^x[38];
	y[5]=x[374]^x[367]^x[352]^x[336]^x[325]^x[315]^x[314]^x[305]^x[304]^x[303]^x[302]^x[294]^x[293]^x[291]^x[251]^x[245]^x[239]^x[234]^x[229]^x[228]^x[214]^x[192]^x[176]^x[165]^x[139]^x[128]^x[101]^x[91]^x[79]^x[74]^x[73]^x[69]^x[67]^x[60]^x[49]^x[37];
	y[4]=x[373]^x[366]^x[362]^x[335]^x[324]^x[314]^x[313]^x[304]^x[303]^x[302]^x[301]^x[293]^x[292]^x[290]^x[250]^x[244]^x[238]^x[233]^x[228]^x[227]^x[213]^x[202]^x[175]^x[164]^x[138]^x[100]^x[90]^x[78]^x[73]^x[72]^x[68]^x[66]^x[59]^x[48]^x[36];
	y[3]=x[372]^x[365]^x[361]^x[334]^x[323]^x[313]^x[312]^x[303]^x[302]^x[301]^x[300]^x[292]^x[291]^x[289]^x[249]^x[243]^x[237]^x[232]^x[227]^x[226]^x[212]^x[201]^x[174]^x[163]^x[137]^x[99]^x[89]^x[77]^x[72]^x[71]^x[67]^x[65]^x[58]^x[47]^x[35];
	y[2]=x[371]^x[364]^x[360]^x[333]^x[322]^x[312]^x[311]^x[302]^x[301]^x[300]^x[299]^x[291]^x[290]^x[288]^x[248]^x[242]^x[236]^x[231]^x[226]^x[225]^x[211]^x[200]^x[173]^x[162]^x[136]^x[98]^x[88]^x[76]^x[71]^x[70]^x[66]^x[64]^x[57]^x[46]^x[34];
	y[1]=x[370]^x[363]^x[359]^x[332]^x[321]^x[311]^x[310]^x[301]^x[300]^x[299]^x[290]^x[289]^x[247]^x[241]^x[235]^x[230]^x[225]^x[224]^x[210]^x[199]^x[172]^x[161]^x[135]^x[97]^x[87]^x[75]^x[70]^x[69]^x[65]^x[56]^x[45]^x[33];
	y[0]=x[369]^x[363]^x[358]^x[352]^x[331]^x[320]^x[310]^x[300]^x[299]^x[289]^x[288]^x[246]^x[240]^x[229]^x[224]^x[209]^x[198]^x[171]^x[160]^x[134]^x[96]^x[86]^x[69]^x[64]^x[55]^x[44]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint47(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[351]^x[346]^x[341]^x[336]^x[330]^x[325]^x[319]^x[313]^x[309]^x[303]^x[298]^x[292]^x[285]^x[278]^x[276]^x[274]^x[267]^x[266]^x[263]^x[223]^x[221]^x[213]^x[212]^x[211]^x[203]^x[201]^x[199]^x[192]^x[186]^x[176]^x[165]^x[159]^x[149]^x[138]^x[122]^x[110]^x[95]^x[83]^x[63]^x[61]^x[57]^x[55]^x[53]^x[52]^x[47]^x[46]^x[43]^x[40]^x[39]^x[37]^x[34]^x[33]^x[32]^x[31]^x[12]^x[11]^x[1];
	y[30]=x[318]^x[312]^x[308]^x[302]^x[297]^x[291]^x[286]^x[284]^x[277]^x[274]^x[273]^x[266]^x[265]^x[263]^x[262]^x[223]^x[222]^x[220]^x[212]^x[211]^x[210]^x[200]^x[198]^x[158]^x[148]^x[137]^x[94]^x[82]^x[63]^x[62]^x[60]^x[57]^x[56]^x[54]^x[52]^x[46]^x[38]^x[32]^x[30]^x[11]^x[10]^x[0];
	y[29]=x[317]^x[311]^x[307]^x[301]^x[296]^x[290]^x[285]^x[283]^x[276]^x[273]^x[272]^x[265]^x[264]^x[262]^x[261]^x[222]^x[221]^x[219]^x[213]^x[211]^x[210]^x[209]^x[207]^x[202]^x[199]^x[197]^x[196]^x[157]^x[147]^x[136]^x[93]^x[81]^x[62]^x[61]^x[59]^x[56]^x[55]^x[51]^x[45]^x[42]^x[37]^x[31]^x[29]^x[9];
	y[28]=x[316]^x[310]^x[306]^x[300]^x[295]^x[289]^x[284]^x[282]^x[275]^x[272]^x[271]^x[264]^x[263]^x[261]^x[260]^x[221]^x[220]^x[218]^x[212]^x[210]^x[209]^x[208]^x[206]^x[201]^x[198]^x[196]^x[195]^x[156]^x[146]^x[135]^x[92]^x[80]^x[61]^x[60]^x[58]^x[55]^x[54]^x[50]^x[44]^x[41]^x[36]^x[30]^x[28]^x[8];
	y[27]=x[315]^x[309]^x[305]^x[299]^x[294]^x[288]^x[283]^x[281]^x[274]^x[271]^x[270]^x[263]^x[262]^x[260]^x[259]^x[220]^x[219]^x[217]^x[211]^x[209]^x[208]^x[207]^x[205]^x[200]^x[197]^x[195]^x[194]^x[155]^x[145]^x[134]^x[91]^x[79]^x[60]^x[59]^x[57]^x[54]^x[53]^x[49]^x[43]^x[40]^x[35]^x[29]^x[27]^x[7];
	y[26]=x[346]^x[341]^x[335]^x[331]^x[320]^x[319]^x[314]^x[308]^x[304]^x[293]^x[282]^x[280]^x[273]^x[270]^x[269]^x[262]^x[261]^x[259]^x[258]^x[223]^x[222]^x[219]^x[218]^x[217]^x[211]^x[208]^x[207]^x[206]^x[205]^x[196]^x[194]^x[181]^x[171]^x[160]^x[154]^x[144]^x[133]^x[117]^x[116]^x[115]^x[90]^x[78]^x[63]^x[62]^x[59]^x[58]^x[56]^x[53]^x[52]^x[51]^x[50]^x[48]^x[42]^x[34]^x[28]^x[26]^x[6];
	y[25]=x[340]^x[334]^x[318]^x[313]^x[307]^x[303]^x[292]^x[281]^x[279]^x[272]^x[269]^x[268]^x[261]^x[260]^x[258]^x[257]^x[222]^x[221]^x[218]^x[217]^x[216]^x[210]^x[207]^x[206]^x[205]^x[204]^x[195]^x[193]^x[180]^x[153]^x[143]^x[132]^x[127]^x[116]^x[114]^x[106]^x[89]^x[77]^x[62]^x[61]^x[58]^x[57]^x[55]^x[52]^x[51]^x[50]^x[49]^x[47]^x[41]^x[33]^x[27]^x[25]^x[5];
	y[24]=x[339]^x[333]^x[317]^x[312]^x[306]^x[302]^x[291]^x[280]^x[278]^x[271]^x[268]^x[267]^x[260]^x[259]^x[257]^x[256]^x[221]^x[220]^x[217]^x[216]^x[215]^x[209]^x[206]^x[205]^x[204]^x[203]^x[194]^x[192]^x[179]^x[152]^x[142]^x[131]^x[126]^x[115]^x[113]^x[105]^x[88]^x[76]^x[61]^x[60]^x[57]^x[56]^x[54]^x[51]^x[50]^x[49]^x[48]^x[46]^x[40]^x[32]^x[26]^x[24]^x[4];
	y[23]=x[338]^x[332]^x[316]^x[311]^x[305]^x[301]^x[290]^x[279]^x[270]^x[259]^x[258]^x[220]^x[219]^x[216]^x[215]^x[214]^x[213]^x[208]^x[207]^x[205]^x[204]^x[203]^x[202]^x[196]^x[193]^x[178]^x[151]^x[141]^x[130]^x[125]^x[114]^x[112]^x[104]^x[87]^x[75]^x[60]^x[59]^x[56]^x[55]^x[50]^x[49]^x[48]^x[47]^x[45]^x[39]^x[36]^x[25]^x[23]^x[3];
	y[22]=x[337]^x[331]^x[315]^x[310]^x[304]^x[300]^x[289]^x[278]^x[269]^x[258]^x[257]^x[219]^x[218]^x[215]^x[214]^x[213]^x[212]^x[207]^x[206]^x[204]^x[203]^x[202]^x[201]^x[195]^x[192]^x[177]^x[150]^x[140]^x[129]^x[124]^x[113]^x[111]^x[103]^x[86]^x[74]^x[59]^x[58]^x[55]^x[54]^x[49]^x[48]^x[47]^x[46]^x[44]^x[38]^x[35]^x[24]^x[22]^x[2];
	y[21]=x[336]^x[331]^x[320]^x[314]^x[309]^x[303]^x[299]^x[288]^x[268]^x[266]^x[257]^x[256]^x[218]^x[217]^x[214]^x[213]^x[212]^x[211]^x[206]^x[205]^x[203]^x[201]^x[200]^x[194]^x[176]^x[149]^x[139]^x[128]^x[123]^x[112]^x[110]^x[102]^x[85]^x[73]^x[58]^x[57]^x[54]^x[53]^x[48]^x[47]^x[46]^x[45]^x[43]^x[42]^x[37]^x[36]^x[34]^x[23]^x[21]^x[1];
	y[20]=x[351]^x[350]^x[346]^x[329]^x[319]^x[313]^x[308]^x[302]^x[287]^x[286]^x[285]^x[276]^x[274]^x[267]^x[266]^x[256]^x[222]^x[213]^x[212]^x[202]^x[200]^x[186]^x[159]^x[148]^x[122]^x[110]^x[101]^x[84]^x[72]^x[62]^x[56]^x[53]^x[52]^x[50]^x[47]^x[46]^x[44]^x[42]^x[41]^x[36]^x[35]^x[22]^x[20]^x[0];
	y[19]=x[349]^x[339]^x[328]^x[318]^x[312]^x[307]^x[301]^x[287]^x[286]^x[285]^x[284]^x[275]^x[273]^x[265]^x[221]^x[212]^x[211]^x[201]^x[199]^x[158]^x[147]^x[83]^x[71]^x[61]^x[55]^x[52]^x[51]^x[49]^x[46]^x[45]^x[43]^x[41]^x[40]^x[35]^x[34]^x[31]^x[21]^x[19]^x[10];
	y[18]=x[348]^x[338]^x[327]^x[317]^x[311]^x[306]^x[300]^x[286]^x[285]^x[284]^x[283]^x[274]^x[272]^x[264]^x[220]^x[211]^x[210]^x[200]^x[198]^x[157]^x[146]^x[82]^x[70]^x[60]^x[54]^x[51]^x[50]^x[48]^x[45]^x[44]^x[42]^x[40]^x[39]^x[34]^x[33]^x[30]^x[20]^x[18]^x[9];
	y[17]=x[347]^x[337]^x[326]^x[316]^x[310]^x[305]^x[299]^x[285]^x[284]^x[283]^x[282]^x[273]^x[271]^x[263]^x[219]^x[213]^x[210]^x[209]^x[207]^x[202]^x[199]^x[197]^x[196]^x[156]^x[145]^x[107]^x[106]^x[96]^x[81]^x[69]^x[59]^x[50]^x[49]^x[47]^x[44]^x[43]^x[42]^x[41]^x[39]^x[38]^x[33]^x[32]^x[29]^x[19]^x[17]^x[8];
	y[16]=x[346]^x[336]^x[325]^x[315]^x[309]^x[304]^x[298]^x[284]^x[283]^x[282]^x[281]^x[272]^x[270]^x[262]^x[218]^x[212]^x[209]^x[208]^x[206]^x[201]^x[198]^x[196]^x[195]^x[155]^x[144]^x[105]^x[80]^x[68]^x[58]^x[49]^x[48]^x[46]^x[43]^x[42]^x[41]^x[40]^x[38]^x[37]^x[32]^x[28]^x[18]^x[16]^x[7];
	y[15]=x[345]^x[341]^x[330]^x[314]^x[308]^x[303]^x[297]^x[283]^x[282]^x[281]^x[280]^x[271]^x[269]^x[261]^x[217]^x[211]^x[208]^x[207]^x[205]^x[200]^x[197]^x[195]^x[194]^x[181]^x[170]^x[154]^x[143]^x[106]^x[104]^x[79]^x[67]^x[57]^x[48]^x[47]^x[45]^x[42]^x[41]^x[40]^x[39]^x[37]^x[36]^x[27]^x[17]^x[15]^x[6];
	y[14]=x[344]^x[340]^x[329]^x[313]^x[307]^x[302]^x[296]^x[282]^x[281]^x[280]^x[279]^x[270]^x[268]^x[260]^x[216]^x[210]^x[207]^x[206]^x[204]^x[199]^x[196]^x[194]^x[193]^x[180]^x[169]^x[153]^x[142]^x[105]^x[103]^x[78]^x[66]^x[56]^x[47]^x[46]^x[44]^x[41]^x[40]^x[39]^x[38]^x[36]^x[35]^x[26]^x[16]^x[14]^x[5];
	y[13]=x[343]^x[339]^x[328]^x[312]^x[306]^x[301]^x[295]^x[281]^x[280]^x[279]^x[278]^x[269]^x[267]^x[259]^x[215]^x[209]^x[206]^x[205]^x[203]^x[198]^x[195]^x[193]^x[192]^x[179]^x[168]^x[152]^x[141]^x[104]^x[102]^x[77]^x[65]^x[55]^x[46]^x[45]^x[43]^x[40]^x[39]^x[38]^x[37]^x[35]^x[34]^x[25]^x[15]^x[13]^x[4];
	y[12]=x[342]^x[338]^x[327]^x[311]^x[305]^x[300]^x[294]^x[280]^x[279]^x[278]^x[268]^x[258]^x[214]^x[208]^x[205]^x[204]^x[197]^x[194]^x[192]^x[178]^x[167]^x[151]^x[140]^x[103]^x[101]^x[76]^x[64]^x[54]^x[45]^x[44]^x[39]^x[38]^x[37]^x[34]^x[33]^x[24]^x[14]^x[12]^x[3];
	y[11]=x[342]^x[337]^x[331]^x[326]^x[310]^x[304]^x[299]^x[293]^x[279]^x[278]^x[257]^x[256]^x[204]^x[203]^x[193]^x[177]^x[166]^x[150]^x[139]^x[102]^x[101]^x[75]^x[44]^x[43]^x[38]^x[37]^x[33]^x[32]^x[23]^x[13]^x[11]^x[2];
	y[10]=x[336]^x[325]^x[309]^x[303]^x[298]^x[292]^x[278]^x[277]^x[266]^x[256]^x[203]^x[202]^x[192]^x[176]^x[165]^x[149]^x[138]^x[101]^x[74]^x[43]^x[42]^x[37]^x[36]^x[32]^x[22]^x[12]^x[10]^x[1];
	y[9]=x[340]^x[339]^x[329]^x[308]^x[302]^x[297]^x[291]^x[287]^x[286]^x[277]^x[276]^x[275]^x[274]^x[266]^x[265]^x[263]^x[223]^x[201]^x[148]^x[137]^x[73]^x[63]^x[57]^x[51]^x[45]^x[41]^x[39]^x[35]^x[33]^x[21]^x[11]^x[9]^x[0];
	y[8]=x[339]^x[338]^x[328]^x[307]^x[301]^x[296]^x[290]^x[286]^x[285]^x[276]^x[275]^x[274]^x[273]^x[265]^x[264]^x[262]^x[222]^x[200]^x[147]^x[136]^x[72]^x[62]^x[56]^x[50]^x[44]^x[40]^x[38]^x[34]^x[32]^x[31]^x[20]^x[8];
	y[7]=x[338]^x[337]^x[327]^x[306]^x[300]^x[295]^x[289]^x[285]^x[284]^x[275]^x[274]^x[273]^x[272]^x[264]^x[263]^x[261]^x[221]^x[199]^x[146]^x[135]^x[71]^x[61]^x[55]^x[49]^x[43]^x[39]^x[37]^x[33]^x[30]^x[19]^x[7];
	y[6]=x[337]^x[336]^x[326]^x[305]^x[299]^x[294]^x[288]^x[284]^x[283]^x[274]^x[273]^x[272]^x[271]^x[263]^x[262]^x[260]^x[220]^x[198]^x[145]^x[134]^x[70]^x[60]^x[54]^x[48]^x[42]^x[38]^x[36]^x[32]^x[29]^x[18]^x[6];
	y[5]=x[342]^x[335]^x[320]^x[304]^x[293]^x[283]^x[282]^x[273]^x[272]^x[271]^x[270]^x[262]^x[261]^x[259]^x[219]^x[213]^x[207]^x[202]^x[197]^x[196]^x[182]^x[160]^x[144]^x[133]^x[107]^x[96]^x[69]^x[59]^x[47]^x[42]^x[41]^x[37]^x[35]^x[28]^x[17]^x[5];
	y[4]=x[341]^x[334]^x[330]^x[303]^x[292]^x[282]^x[281]^x[272]^x[271]^x[270]^x[269]^x[261]^x[260]^x[258]^x[218]^x[212]^x[206]^x[201]^x[196]^x[195]^x[181]^x[170]^x[143]^x[132]^x[106]^x[68]^x[58]^x[46]^x[41]^x[40]^x[36]^x[34]^x[27]^x[16]^x[4];
	y[3]=x[340]^x[333]^x[329]^x[302]^x[291]^x[281]^x[280]^x[271]^x[270]^x[269]^x[268]^x[260]^x[259]^x[257]^x[217]^x[211]^x[205]^x[200]^x[195]^x[194]^x[180]^x[169]^x[142]^x[131]^x[105]^x[67]^x[57]^x[45]^x[40]^x[39]^x[35]^x[33]^x[26]^x[15]^x[3];
	y[2]=x[339]^x[332]^x[328]^x[301]^x[290]^x[280]^x[279]^x[270]^x[269]^x[268]^x[267]^x[259]^x[258]^x[256]^x[216]^x[210]^x[204]^x[199]^x[194]^x[193]^x[179]^x[168]^x[141]^x[130]^x[104]^x[66]^x[56]^x[44]^x[39]^x[38]^x[34]^x[32]^x[25]^x[14]^x[2];
	y[1]=x[338]^x[331]^x[327]^x[300]^x[289]^x[279]^x[278]^x[269]^x[268]^x[267]^x[258]^x[257]^x[215]^x[209]^x[203]^x[198]^x[193]^x[192]^x[178]^x[167]^x[140]^x[129]^x[103]^x[65]^x[55]^x[43]^x[38]^x[37]^x[33]^x[24]^x[13]^x[1];
	y[0]=x[337]^x[331]^x[326]^x[320]^x[299]^x[288]^x[278]^x[268]^x[267]^x[257]^x[256]^x[214]^x[208]^x[197]^x[192]^x[177]^x[166]^x[139]^x[128]^x[102]^x[64]^x[54]^x[37]^x[32]^x[23]^x[12]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint48(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[375]^x[374]^x[373]^x[363]^x[362]^x[353]^x[319]^x[314]^x[309]^x[304]^x[298]^x[293]^x[287]^x[281]^x[277]^x[271]^x[266]^x[260]^x[253]^x[246]^x[244]^x[242]^x[235]^x[234]^x[231]^x[191]^x[189]^x[181]^x[180]^x[179]^x[171]^x[169]^x[167]^x[160]^x[159]^x[154]^x[153]^x[144]^x[140]^x[139]^x[134]^x[129]^x[127]^x[117]^x[106]^x[90]^x[78]^x[63]^x[51]^x[31]^x[29]^x[25]^x[23]^x[21]^x[20]^x[15]^x[14]^x[11]^x[8]^x[7]^x[5]^x[2]^x[1]^x[0];
	y[30]=x[382]^x[374]^x[373]^x[372]^x[362]^x[361]^x[352]^x[286]^x[280]^x[276]^x[270]^x[265]^x[259]^x[254]^x[252]^x[245]^x[242]^x[241]^x[234]^x[233]^x[231]^x[230]^x[191]^x[190]^x[188]^x[180]^x[179]^x[178]^x[168]^x[166]^x[158]^x[152]^x[139]^x[138]^x[133]^x[132]^x[128]^x[126]^x[116]^x[105]^x[62]^x[50]^x[31]^x[30]^x[28]^x[25]^x[24]^x[22]^x[20]^x[14]^x[6]^x[0];
	y[29]=x[383]^x[381]^x[373]^x[372]^x[371]^x[362]^x[361]^x[360]^x[285]^x[279]^x[275]^x[269]^x[264]^x[258]^x[253]^x[251]^x[244]^x[241]^x[240]^x[233]^x[232]^x[230]^x[229]^x[190]^x[189]^x[187]^x[181]^x[179]^x[178]^x[177]^x[175]^x[170]^x[167]^x[165]^x[164]^x[159]^x[157]^x[153]^x[151]^x[137]^x[131]^x[125]^x[115]^x[104]^x[61]^x[49]^x[30]^x[29]^x[27]^x[24]^x[23]^x[19]^x[13]^x[10]^x[5];
	y[28]=x[382]^x[380]^x[372]^x[371]^x[370]^x[361]^x[360]^x[359]^x[284]^x[278]^x[274]^x[268]^x[263]^x[257]^x[252]^x[250]^x[243]^x[240]^x[239]^x[232]^x[231]^x[229]^x[228]^x[189]^x[188]^x[186]^x[180]^x[178]^x[177]^x[176]^x[174]^x[169]^x[166]^x[164]^x[163]^x[158]^x[156]^x[152]^x[150]^x[136]^x[130]^x[124]^x[114]^x[103]^x[60]^x[48]^x[29]^x[28]^x[26]^x[23]^x[22]^x[18]^x[12]^x[9]^x[4];
	y[27]=x[381]^x[379]^x[371]^x[370]^x[369]^x[360]^x[359]^x[358]^x[283]^x[277]^x[273]^x[267]^x[262]^x[256]^x[251]^x[249]^x[242]^x[239]^x[238]^x[231]^x[230]^x[228]^x[227]^x[188]^x[187]^x[185]^x[179]^x[177]^x[176]^x[175]^x[173]^x[168]^x[165]^x[163]^x[162]^x[157]^x[155]^x[151]^x[149]^x[135]^x[129]^x[123]^x[113]^x[102]^x[59]^x[47]^x[28]^x[27]^x[25]^x[22]^x[21]^x[17]^x[11]^x[8]^x[3];
	y[26]=x[380]^x[378]^x[370]^x[369]^x[368]^x[359]^x[358]^x[357]^x[314]^x[309]^x[303]^x[299]^x[288]^x[287]^x[282]^x[276]^x[272]^x[261]^x[250]^x[248]^x[241]^x[238]^x[237]^x[230]^x[229]^x[227]^x[226]^x[191]^x[190]^x[187]^x[186]^x[185]^x[179]^x[176]^x[175]^x[174]^x[173]^x[164]^x[162]^x[156]^x[154]^x[150]^x[149]^x[148]^x[139]^x[134]^x[122]^x[112]^x[101]^x[85]^x[84]^x[83]^x[58]^x[46]^x[31]^x[30]^x[27]^x[26]^x[24]^x[21]^x[20]^x[19]^x[18]^x[16]^x[10]^x[2];
	y[25]=x[379]^x[377]^x[369]^x[368]^x[367]^x[358]^x[357]^x[356]^x[308]^x[302]^x[286]^x[281]^x[275]^x[271]^x[260]^x[249]^x[247]^x[240]^x[237]^x[236]^x[229]^x[228]^x[226]^x[225]^x[190]^x[189]^x[186]^x[185]^x[184]^x[178]^x[175]^x[174]^x[173]^x[172]^x[163]^x[161]^x[155]^x[153]^x[149]^x[148]^x[147]^x[133]^x[121]^x[111]^x[100]^x[95]^x[84]^x[82]^x[74]^x[57]^x[45]^x[30]^x[29]^x[26]^x[25]^x[23]^x[20]^x[19]^x[18]^x[17]^x[15]^x[9]^x[1];
	y[24]=x[378]^x[376]^x[368]^x[367]^x[366]^x[357]^x[356]^x[355]^x[307]^x[301]^x[285]^x[280]^x[274]^x[270]^x[259]^x[248]^x[246]^x[239]^x[236]^x[235]^x[228]^x[227]^x[225]^x[224]^x[189]^x[188]^x[185]^x[184]^x[183]^x[177]^x[174]^x[173]^x[172]^x[171]^x[162]^x[160]^x[154]^x[152]^x[148]^x[147]^x[146]^x[132]^x[120]^x[110]^x[99]^x[94]^x[83]^x[81]^x[73]^x[56]^x[44]^x[29]^x[28]^x[25]^x[24]^x[22]^x[19]^x[18]^x[17]^x[16]^x[14]^x[8]^x[0];
	y[23]=x[377]^x[375]^x[367]^x[366]^x[365]^x[356]^x[355]^x[354]^x[306]^x[300]^x[284]^x[279]^x[273]^x[269]^x[258]^x[247]^x[238]^x[227]^x[226]^x[188]^x[187]^x[184]^x[183]^x[182]^x[181]^x[176]^x[175]^x[173]^x[172]^x[171]^x[170]^x[164]^x[161]^x[153]^x[151]^x[147]^x[146]^x[145]^x[131]^x[119]^x[109]^x[98]^x[93]^x[82]^x[80]^x[72]^x[55]^x[43]^x[28]^x[27]^x[24]^x[23]^x[18]^x[17]^x[16]^x[15]^x[13]^x[7]^x[4];
	y[22]=x[376]^x[374]^x[366]^x[365]^x[364]^x[355]^x[354]^x[353]^x[305]^x[299]^x[283]^x[278]^x[272]^x[268]^x[257]^x[246]^x[237]^x[226]^x[225]^x[187]^x[186]^x[183]^x[182]^x[181]^x[180]^x[175]^x[174]^x[172]^x[171]^x[170]^x[169]^x[163]^x[160]^x[152]^x[150]^x[146]^x[145]^x[144]^x[130]^x[118]^x[108]^x[97]^x[92]^x[81]^x[79]^x[71]^x[54]^x[42]^x[27]^x[26]^x[23]^x[22]^x[17]^x[16]^x[15]^x[14]^x[12]^x[6]^x[3];
	y[21]=x[375]^x[373]^x[365]^x[364]^x[363]^x[354]^x[353]^x[352]^x[304]^x[299]^x[288]^x[282]^x[277]^x[271]^x[267]^x[256]^x[236]^x[234]^x[225]^x[224]^x[186]^x[185]^x[182]^x[181]^x[180]^x[179]^x[174]^x[173]^x[171]^x[169]^x[168]^x[162]^x[151]^x[149]^x[145]^x[144]^x[143]^x[129]^x[117]^x[107]^x[96]^x[91]^x[80]^x[78]^x[70]^x[53]^x[41]^x[26]^x[25]^x[22]^x[21]^x[16]^x[15]^x[14]^x[13]^x[11]^x[10]^x[5]^x[4]^x[2];
	y[20]=x[383]^x[374]^x[372]^x[364]^x[363]^x[353]^x[352]^x[319]^x[318]^x[314]^x[297]^x[287]^x[281]^x[276]^x[270]^x[255]^x[254]^x[253]^x[244]^x[242]^x[235]^x[234]^x[224]^x[190]^x[181]^x[180]^x[170]^x[168]^x[154]^x[150]^x[148]^x[144]^x[142]^x[128]^x[127]^x[116]^x[90]^x[78]^x[69]^x[52]^x[40]^x[30]^x[24]^x[21]^x[20]^x[18]^x[15]^x[14]^x[12]^x[10]^x[9]^x[4]^x[3];
	y[19]=x[383]^x[382]^x[373]^x[371]^x[363]^x[352]^x[317]^x[307]^x[296]^x[286]^x[280]^x[275]^x[269]^x[255]^x[254]^x[253]^x[252]^x[243]^x[241]^x[233]^x[189]^x[180]^x[179]^x[169]^x[167]^x[159]^x[153]^x[149]^x[147]^x[143]^x[141]^x[138]^x[132]^x[126]^x[115]^x[51]^x[39]^x[29]^x[23]^x[20]^x[19]^x[17]^x[14]^x[13]^x[11]^x[9]^x[8]^x[3]^x[2];
	y[18]=x[383]^x[382]^x[381]^x[372]^x[370]^x[316]^x[306]^x[295]^x[285]^x[279]^x[274]^x[268]^x[254]^x[253]^x[252]^x[251]^x[242]^x[240]^x[232]^x[188]^x[179]^x[178]^x[168]^x[166]^x[158]^x[152]^x[148]^x[146]^x[142]^x[140]^x[137]^x[131]^x[125]^x[114]^x[50]^x[38]^x[28]^x[22]^x[19]^x[18]^x[16]^x[13]^x[12]^x[10]^x[8]^x[7]^x[2]^x[1];
	y[17]=x[382]^x[381]^x[380]^x[371]^x[369]^x[315]^x[305]^x[294]^x[284]^x[278]^x[273]^x[267]^x[253]^x[252]^x[251]^x[250]^x[241]^x[239]^x[231]^x[187]^x[181]^x[178]^x[177]^x[175]^x[170]^x[167]^x[165]^x[164]^x[157]^x[151]^x[147]^x[145]^x[141]^x[139]^x[136]^x[130]^x[124]^x[113]^x[75]^x[74]^x[64]^x[49]^x[37]^x[27]^x[18]^x[17]^x[15]^x[12]^x[11]^x[10]^x[9]^x[7]^x[6]^x[1]^x[0];
	y[16]=x[381]^x[380]^x[379]^x[370]^x[368]^x[314]^x[304]^x[293]^x[283]^x[277]^x[272]^x[266]^x[252]^x[251]^x[250]^x[249]^x[240]^x[238]^x[230]^x[186]^x[180]^x[177]^x[176]^x[174]^x[169]^x[166]^x[164]^x[163]^x[156]^x[150]^x[146]^x[144]^x[140]^x[138]^x[135]^x[129]^x[123]^x[112]^x[73]^x[48]^x[36]^x[26]^x[17]^x[16]^x[14]^x[11]^x[10]^x[9]^x[8]^x[6]^x[5]^x[0];
	y[15]=x[380]^x[379]^x[378]^x[369]^x[367]^x[313]^x[309]^x[298]^x[282]^x[276]^x[271]^x[265]^x[251]^x[250]^x[249]^x[248]^x[239]^x[237]^x[229]^x[185]^x[179]^x[176]^x[175]^x[173]^x[168]^x[165]^x[163]^x[162]^x[155]^x[145]^x[143]^x[139]^x[138]^x[137]^x[134]^x[128]^x[122]^x[111]^x[74]^x[72]^x[47]^x[35]^x[25]^x[16]^x[15]^x[13]^x[10]^x[9]^x[8]^x[7]^x[5]^x[4];
	y[14]=x[379]^x[378]^x[377]^x[368]^x[366]^x[312]^x[308]^x[297]^x[281]^x[275]^x[270]^x[264]^x[250]^x[249]^x[248]^x[247]^x[238]^x[236]^x[228]^x[184]^x[178]^x[175]^x[174]^x[172]^x[167]^x[164]^x[162]^x[161]^x[154]^x[144]^x[142]^x[138]^x[137]^x[136]^x[133]^x[121]^x[110]^x[73]^x[71]^x[46]^x[34]^x[24]^x[15]^x[14]^x[12]^x[9]^x[8]^x[7]^x[6]^x[4]^x[3];
	y[13]=x[378]^x[377]^x[376]^x[367]^x[365]^x[311]^x[307]^x[296]^x[280]^x[274]^x[269]^x[263]^x[249]^x[248]^x[247]^x[246]^x[237]^x[235]^x[227]^x[183]^x[177]^x[174]^x[173]^x[171]^x[166]^x[163]^x[161]^x[160]^x[153]^x[143]^x[141]^x[137]^x[136]^x[135]^x[132]^x[120]^x[109]^x[72]^x[70]^x[45]^x[33]^x[23]^x[14]^x[13]^x[11]^x[8]^x[7]^x[6]^x[5]^x[3]^x[2];
	y[12]=x[377]^x[376]^x[375]^x[366]^x[364]^x[310]^x[306]^x[295]^x[279]^x[273]^x[268]^x[262]^x[248]^x[247]^x[246]^x[236]^x[226]^x[182]^x[176]^x[173]^x[172]^x[165]^x[162]^x[160]^x[152]^x[142]^x[140]^x[136]^x[135]^x[134]^x[131]^x[119]^x[108]^x[71]^x[69]^x[44]^x[32]^x[22]^x[13]^x[12]^x[7]^x[6]^x[5]^x[2]^x[1];
	y[11]=x[376]^x[375]^x[374]^x[365]^x[363]^x[310]^x[305]^x[299]^x[294]^x[278]^x[272]^x[267]^x[261]^x[247]^x[246]^x[225]^x[224]^x[172]^x[171]^x[161]^x[151]^x[141]^x[139]^x[135]^x[134]^x[133]^x[130]^x[118]^x[107]^x[70]^x[69]^x[43]^x[12]^x[11]^x[6]^x[5]^x[1]^x[0];
	y[10]=x[375]^x[374]^x[373]^x[364]^x[362]^x[304]^x[293]^x[277]^x[271]^x[266]^x[260]^x[246]^x[245]^x[234]^x[224]^x[171]^x[170]^x[160]^x[150]^x[140]^x[138]^x[134]^x[133]^x[132]^x[129]^x[117]^x[106]^x[69]^x[42]^x[11]^x[10]^x[5]^x[4]^x[0];
	y[9]=x[374]^x[373]^x[372]^x[363]^x[361]^x[308]^x[307]^x[297]^x[276]^x[270]^x[265]^x[259]^x[255]^x[254]^x[245]^x[244]^x[243]^x[242]^x[234]^x[233]^x[231]^x[191]^x[169]^x[149]^x[143]^x[139]^x[137]^x[133]^x[131]^x[128]^x[116]^x[105]^x[41]^x[31]^x[25]^x[19]^x[13]^x[9]^x[7]^x[3]^x[1];
	y[8]=x[373]^x[372]^x[371]^x[362]^x[360]^x[307]^x[306]^x[296]^x[275]^x[269]^x[264]^x[258]^x[254]^x[253]^x[244]^x[243]^x[242]^x[241]^x[233]^x[232]^x[230]^x[190]^x[168]^x[159]^x[153]^x[148]^x[142]^x[136]^x[130]^x[115]^x[104]^x[40]^x[30]^x[24]^x[18]^x[12]^x[8]^x[6]^x[2]^x[0];
	y[7]=x[372]^x[371]^x[370]^x[361]^x[359]^x[306]^x[305]^x[295]^x[274]^x[268]^x[263]^x[257]^x[253]^x[252]^x[243]^x[242]^x[241]^x[240]^x[232]^x[231]^x[229]^x[189]^x[167]^x[158]^x[152]^x[147]^x[141]^x[135]^x[129]^x[114]^x[103]^x[39]^x[29]^x[23]^x[17]^x[11]^x[7]^x[5]^x[1];
	y[6]=x[371]^x[370]^x[369]^x[360]^x[358]^x[305]^x[304]^x[294]^x[273]^x[267]^x[262]^x[256]^x[252]^x[251]^x[242]^x[241]^x[240]^x[239]^x[231]^x[230]^x[228]^x[188]^x[166]^x[157]^x[151]^x[146]^x[140]^x[134]^x[128]^x[113]^x[102]^x[38]^x[28]^x[22]^x[16]^x[10]^x[6]^x[4]^x[0];
	y[5]=x[370]^x[369]^x[368]^x[359]^x[357]^x[310]^x[303]^x[288]^x[272]^x[261]^x[251]^x[250]^x[241]^x[240]^x[239]^x[238]^x[230]^x[229]^x[227]^x[187]^x[181]^x[175]^x[170]^x[165]^x[164]^x[156]^x[145]^x[139]^x[133]^x[128]^x[112]^x[101]^x[75]^x[64]^x[37]^x[27]^x[15]^x[10]^x[9]^x[5]^x[3];
	y[4]=x[369]^x[368]^x[367]^x[358]^x[356]^x[309]^x[302]^x[298]^x[271]^x[260]^x[250]^x[249]^x[240]^x[239]^x[238]^x[237]^x[229]^x[228]^x[226]^x[186]^x[180]^x[174]^x[169]^x[164]^x[163]^x[155]^x[144]^x[132]^x[111]^x[100]^x[74]^x[36]^x[26]^x[14]^x[9]^x[8]^x[4]^x[2];
	y[3]=x[368]^x[367]^x[366]^x[357]^x[355]^x[308]^x[301]^x[297]^x[270]^x[259]^x[249]^x[248]^x[239]^x[238]^x[237]^x[236]^x[228]^x[227]^x[225]^x[185]^x[179]^x[173]^x[168]^x[163]^x[162]^x[154]^x[143]^x[131]^x[110]^x[99]^x[73]^x[35]^x[25]^x[13]^x[8]^x[7]^x[3]^x[1];
	y[2]=x[367]^x[366]^x[365]^x[356]^x[354]^x[307]^x[300]^x[296]^x[269]^x[258]^x[248]^x[247]^x[238]^x[237]^x[236]^x[235]^x[227]^x[226]^x[224]^x[184]^x[178]^x[172]^x[167]^x[162]^x[161]^x[153]^x[142]^x[130]^x[109]^x[98]^x[72]^x[34]^x[24]^x[12]^x[7]^x[6]^x[2]^x[0];
	y[1]=x[366]^x[365]^x[364]^x[355]^x[353]^x[306]^x[299]^x[295]^x[268]^x[257]^x[247]^x[246]^x[237]^x[236]^x[235]^x[226]^x[225]^x[183]^x[177]^x[171]^x[166]^x[161]^x[160]^x[152]^x[141]^x[129]^x[108]^x[97]^x[71]^x[33]^x[23]^x[11]^x[6]^x[5]^x[1];
	y[0]=x[365]^x[364]^x[363]^x[354]^x[352]^x[305]^x[299]^x[294]^x[288]^x[267]^x[256]^x[246]^x[236]^x[235]^x[225]^x[224]^x[182]^x[176]^x[165]^x[160]^x[151]^x[140]^x[128]^x[107]^x[96]^x[70]^x[32]^x[22]^x[5]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint49(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[381]^x[378]^x[375]^x[374]^x[372]^x[370]^x[368]^x[366]^x[364]^x[363]^x[362]^x[359]^x[357]^x[356]^x[353]^x[351]^x[343]^x[342]^x[341]^x[331]^x[330]^x[321]^x[287]^x[282]^x[277]^x[272]^x[266]^x[261]^x[255]^x[249]^x[245]^x[239]^x[234]^x[228]^x[221]^x[214]^x[212]^x[210]^x[203]^x[202]^x[199]^x[145]^x[127]^x[122]^x[121]^x[112]^x[108]^x[107]^x[102]^x[97]^x[95]^x[85]^x[74]^x[58]^x[46]^x[31]^x[19];
	y[30]=x[382]^x[380]^x[376]^x[374]^x[373]^x[370]^x[369]^x[367]^x[364]^x[363]^x[362]^x[361]^x[359]^x[358]^x[356]^x[355]^x[353]^x[352]^x[350]^x[342]^x[341]^x[340]^x[330]^x[329]^x[320]^x[254]^x[248]^x[244]^x[238]^x[233]^x[227]^x[222]^x[220]^x[213]^x[210]^x[209]^x[202]^x[201]^x[199]^x[198]^x[144]^x[126]^x[120]^x[107]^x[106]^x[101]^x[100]^x[96]^x[94]^x[84]^x[73]^x[30]^x[18];
	y[29]=x[381]^x[379]^x[375]^x[373]^x[372]^x[369]^x[368]^x[366]^x[362]^x[361]^x[360]^x[358]^x[357]^x[355]^x[354]^x[351]^x[349]^x[341]^x[340]^x[339]^x[330]^x[329]^x[328]^x[253]^x[247]^x[243]^x[237]^x[232]^x[226]^x[221]^x[219]^x[212]^x[209]^x[208]^x[201]^x[200]^x[198]^x[197]^x[143]^x[127]^x[125]^x[121]^x[119]^x[105]^x[99]^x[93]^x[83]^x[72]^x[29]^x[17];
	y[28]=x[380]^x[378]^x[374]^x[372]^x[371]^x[368]^x[367]^x[365]^x[361]^x[360]^x[359]^x[357]^x[356]^x[354]^x[353]^x[350]^x[348]^x[340]^x[339]^x[338]^x[329]^x[328]^x[327]^x[252]^x[246]^x[242]^x[236]^x[231]^x[225]^x[220]^x[218]^x[211]^x[208]^x[207]^x[200]^x[199]^x[197]^x[196]^x[142]^x[126]^x[124]^x[120]^x[118]^x[104]^x[98]^x[92]^x[82]^x[71]^x[28]^x[16];
	y[27]=x[379]^x[377]^x[373]^x[371]^x[370]^x[367]^x[366]^x[364]^x[360]^x[359]^x[358]^x[356]^x[355]^x[353]^x[352]^x[349]^x[347]^x[339]^x[338]^x[337]^x[328]^x[327]^x[326]^x[251]^x[245]^x[241]^x[235]^x[230]^x[224]^x[219]^x[217]^x[210]^x[207]^x[206]^x[199]^x[198]^x[196]^x[195]^x[141]^x[125]^x[123]^x[119]^x[117]^x[103]^x[97]^x[91]^x[81]^x[70]^x[27]^x[15];
	y[26]=x[381]^x[378]^x[376]^x[373]^x[371]^x[370]^x[369]^x[366]^x[365]^x[363]^x[361]^x[358]^x[357]^x[355]^x[354]^x[352]^x[348]^x[346]^x[338]^x[337]^x[336]^x[327]^x[326]^x[325]^x[282]^x[277]^x[271]^x[267]^x[256]^x[255]^x[250]^x[244]^x[240]^x[229]^x[218]^x[216]^x[209]^x[206]^x[205]^x[198]^x[197]^x[195]^x[194]^x[140]^x[124]^x[122]^x[118]^x[117]^x[116]^x[107]^x[102]^x[90]^x[80]^x[69]^x[53]^x[52]^x[51]^x[26]^x[14];
	y[25]=x[383]^x[380]^x[377]^x[375]^x[372]^x[370]^x[369]^x[368]^x[365]^x[364]^x[360]^x[357]^x[356]^x[354]^x[353]^x[347]^x[345]^x[337]^x[336]^x[335]^x[326]^x[325]^x[324]^x[276]^x[270]^x[254]^x[249]^x[243]^x[239]^x[228]^x[217]^x[215]^x[208]^x[205]^x[204]^x[197]^x[196]^x[194]^x[193]^x[139]^x[123]^x[121]^x[117]^x[116]^x[115]^x[101]^x[89]^x[79]^x[68]^x[63]^x[52]^x[50]^x[42]^x[25]^x[13];
	y[24]=x[382]^x[379]^x[376]^x[374]^x[371]^x[369]^x[368]^x[367]^x[364]^x[363]^x[359]^x[356]^x[355]^x[353]^x[352]^x[346]^x[344]^x[336]^x[335]^x[334]^x[325]^x[324]^x[323]^x[275]^x[269]^x[253]^x[248]^x[242]^x[238]^x[227]^x[216]^x[214]^x[207]^x[204]^x[203]^x[196]^x[195]^x[193]^x[192]^x[138]^x[122]^x[120]^x[116]^x[115]^x[114]^x[100]^x[88]^x[78]^x[67]^x[62]^x[51]^x[49]^x[41]^x[24]^x[12];
	y[23]=x[381]^x[378]^x[375]^x[370]^x[368]^x[366]^x[358]^x[356]^x[355]^x[354]^x[345]^x[343]^x[335]^x[334]^x[333]^x[324]^x[323]^x[322]^x[274]^x[268]^x[252]^x[247]^x[241]^x[237]^x[226]^x[215]^x[206]^x[195]^x[194]^x[137]^x[121]^x[119]^x[115]^x[114]^x[113]^x[99]^x[87]^x[77]^x[66]^x[61]^x[50]^x[48]^x[40]^x[23]^x[11];
	y[22]=x[380]^x[377]^x[374]^x[369]^x[367]^x[365]^x[357]^x[355]^x[354]^x[353]^x[344]^x[342]^x[334]^x[333]^x[332]^x[323]^x[322]^x[321]^x[273]^x[267]^x[251]^x[246]^x[240]^x[236]^x[225]^x[214]^x[205]^x[194]^x[193]^x[136]^x[120]^x[118]^x[114]^x[113]^x[112]^x[98]^x[86]^x[76]^x[65]^x[60]^x[49]^x[47]^x[39]^x[22]^x[10];
	y[21]=x[379]^x[376]^x[368]^x[367]^x[366]^x[364]^x[362]^x[354]^x[353]^x[352]^x[343]^x[341]^x[333]^x[332]^x[331]^x[322]^x[321]^x[320]^x[272]^x[267]^x[256]^x[250]^x[245]^x[239]^x[235]^x[224]^x[204]^x[202]^x[193]^x[192]^x[135]^x[119]^x[117]^x[113]^x[112]^x[111]^x[97]^x[85]^x[75]^x[64]^x[59]^x[48]^x[46]^x[38]^x[21]^x[9];
	y[20]=x[383]^x[382]^x[381]^x[378]^x[377]^x[376]^x[375]^x[372]^x[370]^x[366]^x[364]^x[363]^x[362]^x[356]^x[352]^x[351]^x[342]^x[340]^x[332]^x[331]^x[321]^x[320]^x[287]^x[286]^x[282]^x[265]^x[255]^x[249]^x[244]^x[238]^x[223]^x[222]^x[221]^x[212]^x[210]^x[203]^x[202]^x[192]^x[134]^x[122]^x[118]^x[116]^x[112]^x[110]^x[96]^x[95]^x[84]^x[58]^x[46]^x[37]^x[20]^x[8];
	y[19]=x[383]^x[382]^x[381]^x[380]^x[377]^x[376]^x[375]^x[374]^x[371]^x[369]^x[365]^x[363]^x[361]^x[355]^x[351]^x[350]^x[341]^x[339]^x[331]^x[320]^x[285]^x[275]^x[264]^x[254]^x[248]^x[243]^x[237]^x[223]^x[222]^x[221]^x[220]^x[211]^x[209]^x[201]^x[133]^x[127]^x[121]^x[117]^x[115]^x[111]^x[109]^x[106]^x[100]^x[94]^x[83]^x[19]^x[7];
	y[18]=x[382]^x[381]^x[380]^x[379]^x[376]^x[375]^x[374]^x[373]^x[370]^x[368]^x[364]^x[362]^x[360]^x[354]^x[351]^x[350]^x[349]^x[340]^x[338]^x[284]^x[274]^x[263]^x[253]^x[247]^x[242]^x[236]^x[222]^x[221]^x[220]^x[219]^x[210]^x[208]^x[200]^x[132]^x[126]^x[120]^x[116]^x[114]^x[110]^x[108]^x[105]^x[99]^x[93]^x[82]^x[18]^x[6];
	y[17]=x[381]^x[380]^x[379]^x[378]^x[375]^x[374]^x[373]^x[372]^x[369]^x[367]^x[362]^x[361]^x[359]^x[353]^x[352]^x[350]^x[349]^x[348]^x[339]^x[337]^x[283]^x[273]^x[262]^x[252]^x[246]^x[241]^x[235]^x[221]^x[220]^x[219]^x[218]^x[209]^x[207]^x[199]^x[131]^x[125]^x[119]^x[115]^x[113]^x[109]^x[107]^x[104]^x[98]^x[92]^x[81]^x[43]^x[42]^x[32]^x[17]^x[5];
	y[16]=x[380]^x[379]^x[378]^x[377]^x[374]^x[373]^x[372]^x[371]^x[368]^x[366]^x[362]^x[361]^x[360]^x[358]^x[352]^x[349]^x[348]^x[347]^x[338]^x[336]^x[282]^x[272]^x[261]^x[251]^x[245]^x[240]^x[234]^x[220]^x[219]^x[218]^x[217]^x[208]^x[206]^x[198]^x[130]^x[124]^x[118]^x[114]^x[112]^x[108]^x[106]^x[103]^x[97]^x[91]^x[80]^x[41]^x[16]^x[4];
	y[15]=x[379]^x[378]^x[377]^x[376]^x[373]^x[372]^x[371]^x[370]^x[367]^x[365]^x[362]^x[361]^x[360]^x[359]^x[357]^x[348]^x[347]^x[346]^x[337]^x[335]^x[281]^x[277]^x[266]^x[250]^x[244]^x[239]^x[233]^x[219]^x[218]^x[217]^x[216]^x[207]^x[205]^x[197]^x[129]^x[123]^x[113]^x[111]^x[107]^x[106]^x[105]^x[102]^x[96]^x[90]^x[79]^x[42]^x[40]^x[15]^x[3];
	y[14]=x[378]^x[377]^x[376]^x[375]^x[372]^x[371]^x[370]^x[369]^x[366]^x[364]^x[361]^x[360]^x[359]^x[358]^x[356]^x[347]^x[346]^x[345]^x[336]^x[334]^x[280]^x[276]^x[265]^x[249]^x[243]^x[238]^x[232]^x[218]^x[217]^x[216]^x[215]^x[206]^x[204]^x[196]^x[128]^x[122]^x[112]^x[110]^x[106]^x[105]^x[104]^x[101]^x[89]^x[78]^x[41]^x[39]^x[14]^x[2];
	y[13]=x[377]^x[376]^x[375]^x[374]^x[371]^x[370]^x[369]^x[368]^x[365]^x[363]^x[360]^x[359]^x[358]^x[357]^x[355]^x[346]^x[345]^x[344]^x[335]^x[333]^x[279]^x[275]^x[264]^x[248]^x[242]^x[237]^x[231]^x[217]^x[216]^x[215]^x[214]^x[205]^x[203]^x[195]^x[121]^x[111]^x[109]^x[105]^x[104]^x[103]^x[100]^x[88]^x[77]^x[40]^x[38]^x[13]^x[1];
	y[12]=x[376]^x[375]^x[374]^x[370]^x[369]^x[368]^x[364]^x[359]^x[358]^x[357]^x[354]^x[345]^x[344]^x[343]^x[334]^x[332]^x[278]^x[274]^x[263]^x[247]^x[241]^x[236]^x[230]^x[216]^x[215]^x[214]^x[204]^x[194]^x[120]^x[110]^x[108]^x[104]^x[103]^x[102]^x[99]^x[87]^x[76]^x[39]^x[37]^x[12]^x[0];
	y[11]=x[375]^x[374]^x[369]^x[368]^x[358]^x[357]^x[353]^x[352]^x[344]^x[343]^x[342]^x[333]^x[331]^x[278]^x[273]^x[267]^x[262]^x[246]^x[240]^x[235]^x[229]^x[215]^x[214]^x[193]^x[192]^x[119]^x[109]^x[107]^x[103]^x[102]^x[101]^x[98]^x[86]^x[75]^x[38]^x[37]^x[11];
	y[10]=x[374]^x[373]^x[368]^x[367]^x[362]^x[357]^x[356]^x[352]^x[343]^x[342]^x[341]^x[332]^x[330]^x[272]^x[261]^x[245]^x[239]^x[234]^x[228]^x[214]^x[213]^x[202]^x[192]^x[118]^x[108]^x[106]^x[102]^x[101]^x[100]^x[97]^x[85]^x[74]^x[37]^x[10];
	y[9]=x[383]^x[382]^x[377]^x[376]^x[373]^x[372]^x[371]^x[370]^x[367]^x[366]^x[365]^x[364]^x[362]^x[361]^x[359]^x[356]^x[355]^x[353]^x[342]^x[341]^x[340]^x[331]^x[329]^x[276]^x[275]^x[265]^x[244]^x[238]^x[233]^x[227]^x[223]^x[222]^x[213]^x[212]^x[211]^x[210]^x[202]^x[201]^x[199]^x[117]^x[111]^x[107]^x[105]^x[101]^x[99]^x[96]^x[84]^x[73]^x[9];
	y[8]=x[382]^x[381]^x[376]^x[375]^x[372]^x[371]^x[370]^x[369]^x[366]^x[365]^x[364]^x[363]^x[361]^x[360]^x[358]^x[355]^x[354]^x[352]^x[341]^x[340]^x[339]^x[330]^x[328]^x[275]^x[274]^x[264]^x[243]^x[237]^x[232]^x[226]^x[222]^x[221]^x[212]^x[211]^x[210]^x[209]^x[201]^x[200]^x[198]^x[127]^x[121]^x[116]^x[110]^x[104]^x[98]^x[83]^x[72]^x[8];
	y[7]=x[381]^x[380]^x[375]^x[374]^x[371]^x[370]^x[369]^x[368]^x[365]^x[364]^x[363]^x[360]^x[359]^x[357]^x[354]^x[353]^x[340]^x[339]^x[338]^x[329]^x[327]^x[274]^x[273]^x[263]^x[242]^x[236]^x[231]^x[225]^x[221]^x[220]^x[211]^x[210]^x[209]^x[208]^x[200]^x[199]^x[197]^x[126]^x[120]^x[115]^x[109]^x[103]^x[97]^x[82]^x[71]^x[7];
	y[6]=x[380]^x[379]^x[374]^x[373]^x[370]^x[369]^x[368]^x[367]^x[364]^x[363]^x[362]^x[359]^x[358]^x[356]^x[353]^x[352]^x[339]^x[338]^x[337]^x[328]^x[326]^x[273]^x[272]^x[262]^x[241]^x[235]^x[230]^x[224]^x[220]^x[219]^x[210]^x[209]^x[208]^x[207]^x[199]^x[198]^x[196]^x[125]^x[119]^x[114]^x[108]^x[102]^x[96]^x[81]^x[70]^x[6];
	y[5]=x[379]^x[378]^x[373]^x[372]^x[369]^x[368]^x[367]^x[366]^x[362]^x[361]^x[358]^x[357]^x[355]^x[338]^x[337]^x[336]^x[327]^x[325]^x[278]^x[271]^x[256]^x[240]^x[229]^x[219]^x[218]^x[209]^x[208]^x[207]^x[206]^x[198]^x[197]^x[195]^x[124]^x[113]^x[107]^x[101]^x[96]^x[80]^x[69]^x[43]^x[32]^x[5];
	y[4]=x[378]^x[377]^x[372]^x[371]^x[368]^x[367]^x[366]^x[365]^x[361]^x[360]^x[357]^x[356]^x[354]^x[337]^x[336]^x[335]^x[326]^x[324]^x[277]^x[270]^x[266]^x[239]^x[228]^x[218]^x[217]^x[208]^x[207]^x[206]^x[205]^x[197]^x[196]^x[194]^x[123]^x[112]^x[100]^x[79]^x[68]^x[42]^x[4];
	y[3]=x[377]^x[376]^x[371]^x[370]^x[367]^x[366]^x[365]^x[364]^x[360]^x[359]^x[356]^x[355]^x[353]^x[336]^x[335]^x[334]^x[325]^x[323]^x[276]^x[269]^x[265]^x[238]^x[227]^x[217]^x[216]^x[207]^x[206]^x[205]^x[204]^x[196]^x[195]^x[193]^x[122]^x[111]^x[99]^x[78]^x[67]^x[41]^x[3];
	y[2]=x[376]^x[375]^x[370]^x[369]^x[366]^x[365]^x[364]^x[363]^x[359]^x[358]^x[355]^x[354]^x[352]^x[335]^x[334]^x[333]^x[324]^x[322]^x[275]^x[268]^x[264]^x[237]^x[226]^x[216]^x[215]^x[206]^x[205]^x[204]^x[203]^x[195]^x[194]^x[192]^x[121]^x[110]^x[98]^x[77]^x[66]^x[40]^x[2];
	y[1]=x[375]^x[374]^x[369]^x[368]^x[365]^x[364]^x[363]^x[358]^x[357]^x[354]^x[353]^x[334]^x[333]^x[332]^x[323]^x[321]^x[274]^x[267]^x[263]^x[236]^x[225]^x[215]^x[214]^x[205]^x[204]^x[203]^x[194]^x[193]^x[120]^x[109]^x[97]^x[76]^x[65]^x[39]^x[1];
	y[0]=x[374]^x[368]^x[364]^x[363]^x[357]^x[353]^x[352]^x[333]^x[332]^x[331]^x[322]^x[320]^x[273]^x[267]^x[262]^x[256]^x[235]^x[224]^x[214]^x[204]^x[203]^x[193]^x[192]^x[119]^x[108]^x[96]^x[75]^x[64]^x[38]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint50(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[373]^x[371]^x[362]^x[349]^x[346]^x[343]^x[342]^x[340]^x[338]^x[336]^x[334]^x[332]^x[331]^x[330]^x[327]^x[325]^x[324]^x[321]^x[319]^x[311]^x[310]^x[309]^x[299]^x[298]^x[289]^x[255]^x[250]^x[245]^x[240]^x[234]^x[229]^x[223]^x[217]^x[213]^x[207]^x[202]^x[196]^x[189]^x[182]^x[180]^x[178]^x[171]^x[170]^x[167]^x[159]^x[153]^x[147]^x[141]^x[113]^x[95]^x[90]^x[89]^x[80]^x[76]^x[75]^x[70]^x[65]^x[63]^x[53]^x[42]^x[26]^x[14];
	y[30]=x[382]^x[381]^x[372]^x[370]^x[361]^x[350]^x[348]^x[344]^x[342]^x[341]^x[338]^x[337]^x[335]^x[332]^x[331]^x[330]^x[329]^x[327]^x[326]^x[324]^x[323]^x[321]^x[320]^x[318]^x[310]^x[309]^x[308]^x[298]^x[297]^x[288]^x[222]^x[216]^x[212]^x[206]^x[201]^x[195]^x[190]^x[188]^x[181]^x[178]^x[177]^x[170]^x[169]^x[167]^x[166]^x[158]^x[152]^x[146]^x[140]^x[112]^x[94]^x[88]^x[75]^x[74]^x[69]^x[68]^x[64]^x[62]^x[52]^x[41];
	y[29]=x[381]^x[380]^x[371]^x[369]^x[360]^x[349]^x[347]^x[343]^x[341]^x[340]^x[337]^x[336]^x[334]^x[330]^x[329]^x[328]^x[326]^x[325]^x[323]^x[322]^x[319]^x[317]^x[309]^x[308]^x[307]^x[298]^x[297]^x[296]^x[221]^x[215]^x[211]^x[205]^x[200]^x[194]^x[189]^x[187]^x[180]^x[177]^x[176]^x[169]^x[168]^x[166]^x[165]^x[157]^x[151]^x[145]^x[139]^x[111]^x[95]^x[93]^x[89]^x[87]^x[73]^x[67]^x[61]^x[51]^x[40];
	y[28]=x[380]^x[379]^x[370]^x[368]^x[359]^x[348]^x[346]^x[342]^x[340]^x[339]^x[336]^x[335]^x[333]^x[329]^x[328]^x[327]^x[325]^x[324]^x[322]^x[321]^x[318]^x[316]^x[308]^x[307]^x[306]^x[297]^x[296]^x[295]^x[220]^x[214]^x[210]^x[204]^x[199]^x[193]^x[188]^x[186]^x[179]^x[176]^x[175]^x[168]^x[167]^x[165]^x[164]^x[156]^x[150]^x[144]^x[138]^x[110]^x[94]^x[92]^x[88]^x[86]^x[72]^x[66]^x[60]^x[50]^x[39];
	y[27]=x[379]^x[378]^x[369]^x[367]^x[358]^x[347]^x[345]^x[341]^x[339]^x[338]^x[335]^x[334]^x[332]^x[328]^x[327]^x[326]^x[324]^x[323]^x[321]^x[320]^x[317]^x[315]^x[307]^x[306]^x[305]^x[296]^x[295]^x[294]^x[219]^x[213]^x[209]^x[203]^x[198]^x[192]^x[187]^x[185]^x[178]^x[175]^x[174]^x[167]^x[166]^x[164]^x[163]^x[155]^x[149]^x[143]^x[137]^x[109]^x[93]^x[91]^x[87]^x[85]^x[71]^x[65]^x[59]^x[49]^x[38];
	y[26]=x[378]^x[377]^x[368]^x[366]^x[357]^x[349]^x[346]^x[344]^x[341]^x[339]^x[338]^x[337]^x[334]^x[333]^x[331]^x[329]^x[326]^x[325]^x[323]^x[322]^x[320]^x[316]^x[314]^x[306]^x[305]^x[304]^x[295]^x[294]^x[293]^x[250]^x[245]^x[239]^x[235]^x[224]^x[223]^x[218]^x[212]^x[208]^x[197]^x[186]^x[184]^x[177]^x[174]^x[173]^x[166]^x[165]^x[163]^x[162]^x[154]^x[148]^x[142]^x[136]^x[108]^x[92]^x[90]^x[86]^x[85]^x[84]^x[75]^x[70]^x[58]^x[48]^x[37]^x[21]^x[20]^x[19];
	y[25]=x[377]^x[376]^x[367]^x[365]^x[356]^x[351]^x[348]^x[345]^x[343]^x[340]^x[338]^x[337]^x[336]^x[333]^x[332]^x[328]^x[325]^x[324]^x[322]^x[321]^x[315]^x[313]^x[305]^x[304]^x[303]^x[294]^x[293]^x[292]^x[244]^x[238]^x[222]^x[217]^x[211]^x[207]^x[196]^x[185]^x[183]^x[176]^x[173]^x[172]^x[165]^x[164]^x[162]^x[161]^x[153]^x[147]^x[141]^x[135]^x[107]^x[91]^x[89]^x[85]^x[84]^x[83]^x[69]^x[57]^x[47]^x[36]^x[31]^x[20]^x[18]^x[10];
	y[24]=x[376]^x[375]^x[366]^x[364]^x[355]^x[350]^x[347]^x[344]^x[342]^x[339]^x[337]^x[336]^x[335]^x[332]^x[331]^x[327]^x[324]^x[323]^x[321]^x[320]^x[314]^x[312]^x[304]^x[303]^x[302]^x[293]^x[292]^x[291]^x[243]^x[237]^x[221]^x[216]^x[210]^x[206]^x[195]^x[184]^x[182]^x[175]^x[172]^x[171]^x[164]^x[163]^x[161]^x[160]^x[152]^x[146]^x[140]^x[134]^x[106]^x[90]^x[88]^x[84]^x[83]^x[82]^x[68]^x[56]^x[46]^x[35]^x[30]^x[19]^x[17]^x[9];
	y[23]=x[375]^x[374]^x[365]^x[363]^x[354]^x[349]^x[346]^x[343]^x[338]^x[336]^x[334]^x[326]^x[324]^x[323]^x[322]^x[313]^x[311]^x[303]^x[302]^x[301]^x[292]^x[291]^x[290]^x[242]^x[236]^x[220]^x[215]^x[209]^x[205]^x[194]^x[183]^x[174]^x[163]^x[162]^x[151]^x[145]^x[139]^x[133]^x[105]^x[89]^x[87]^x[83]^x[82]^x[81]^x[67]^x[55]^x[45]^x[34]^x[29]^x[18]^x[16]^x[8];
	y[22]=x[374]^x[373]^x[364]^x[362]^x[353]^x[348]^x[345]^x[342]^x[337]^x[335]^x[333]^x[325]^x[323]^x[322]^x[321]^x[312]^x[310]^x[302]^x[301]^x[300]^x[291]^x[290]^x[289]^x[241]^x[235]^x[219]^x[214]^x[208]^x[204]^x[193]^x[182]^x[173]^x[162]^x[161]^x[150]^x[144]^x[138]^x[132]^x[104]^x[88]^x[86]^x[82]^x[81]^x[80]^x[66]^x[54]^x[44]^x[33]^x[28]^x[17]^x[15]^x[7];
	y[21]=x[373]^x[372]^x[363]^x[361]^x[352]^x[347]^x[344]^x[336]^x[335]^x[334]^x[332]^x[330]^x[322]^x[321]^x[320]^x[311]^x[309]^x[301]^x[300]^x[299]^x[290]^x[289]^x[288]^x[240]^x[235]^x[224]^x[218]^x[213]^x[207]^x[203]^x[192]^x[172]^x[170]^x[161]^x[160]^x[149]^x[143]^x[137]^x[131]^x[103]^x[87]^x[85]^x[81]^x[80]^x[79]^x[65]^x[53]^x[43]^x[32]^x[27]^x[16]^x[14]^x[6];
	y[20]=x[383]^x[372]^x[371]^x[360]^x[351]^x[350]^x[349]^x[346]^x[345]^x[344]^x[343]^x[340]^x[338]^x[334]^x[332]^x[331]^x[330]^x[324]^x[320]^x[319]^x[310]^x[308]^x[300]^x[299]^x[289]^x[288]^x[255]^x[254]^x[250]^x[233]^x[223]^x[217]^x[212]^x[206]^x[191]^x[190]^x[189]^x[180]^x[178]^x[171]^x[170]^x[160]^x[148]^x[142]^x[136]^x[130]^x[102]^x[90]^x[86]^x[84]^x[80]^x[78]^x[64]^x[63]^x[52]^x[26]^x[14]^x[5];
	y[19]=x[382]^x[371]^x[370]^x[359]^x[351]^x[350]^x[349]^x[348]^x[345]^x[344]^x[343]^x[342]^x[339]^x[337]^x[333]^x[331]^x[329]^x[323]^x[319]^x[318]^x[309]^x[307]^x[299]^x[288]^x[253]^x[243]^x[232]^x[222]^x[216]^x[211]^x[205]^x[191]^x[190]^x[189]^x[188]^x[179]^x[177]^x[169]^x[147]^x[141]^x[135]^x[129]^x[101]^x[95]^x[89]^x[85]^x[83]^x[79]^x[77]^x[74]^x[68]^x[62]^x[51];
	y[18]=x[381]^x[370]^x[369]^x[358]^x[350]^x[349]^x[348]^x[347]^x[344]^x[343]^x[342]^x[341]^x[338]^x[336]^x[332]^x[330]^x[328]^x[322]^x[319]^x[318]^x[317]^x[308]^x[306]^x[252]^x[242]^x[231]^x[221]^x[215]^x[210]^x[204]^x[190]^x[189]^x[188]^x[187]^x[178]^x[176]^x[168]^x[146]^x[140]^x[134]^x[128]^x[100]^x[94]^x[88]^x[84]^x[82]^x[78]^x[76]^x[73]^x[67]^x[61]^x[50];
	y[17]=x[380]^x[369]^x[368]^x[357]^x[349]^x[348]^x[347]^x[346]^x[343]^x[342]^x[341]^x[340]^x[337]^x[335]^x[330]^x[329]^x[327]^x[321]^x[320]^x[318]^x[317]^x[316]^x[307]^x[305]^x[251]^x[241]^x[230]^x[220]^x[214]^x[209]^x[203]^x[189]^x[188]^x[187]^x[186]^x[177]^x[175]^x[167]^x[145]^x[139]^x[133]^x[99]^x[93]^x[87]^x[83]^x[81]^x[77]^x[75]^x[72]^x[66]^x[60]^x[49]^x[11]^x[10]^x[0];
	y[16]=x[379]^x[368]^x[367]^x[356]^x[348]^x[347]^x[346]^x[345]^x[342]^x[341]^x[340]^x[339]^x[336]^x[334]^x[330]^x[329]^x[328]^x[326]^x[320]^x[317]^x[316]^x[315]^x[306]^x[304]^x[250]^x[240]^x[229]^x[219]^x[213]^x[208]^x[202]^x[188]^x[187]^x[186]^x[185]^x[176]^x[174]^x[166]^x[144]^x[138]^x[132]^x[98]^x[92]^x[86]^x[82]^x[80]^x[76]^x[74]^x[71]^x[65]^x[59]^x[48]^x[9];
	y[15]=x[378]^x[367]^x[366]^x[355]^x[347]^x[346]^x[345]^x[344]^x[341]^x[340]^x[339]^x[338]^x[335]^x[333]^x[330]^x[329]^x[328]^x[327]^x[325]^x[316]^x[315]^x[314]^x[305]^x[303]^x[249]^x[245]^x[234]^x[218]^x[212]^x[207]^x[201]^x[187]^x[186]^x[185]^x[184]^x[175]^x[173]^x[165]^x[143]^x[137]^x[131]^x[97]^x[91]^x[81]^x[79]^x[75]^x[74]^x[73]^x[70]^x[64]^x[58]^x[47]^x[10]^x[8];
	y[14]=x[377]^x[366]^x[365]^x[354]^x[346]^x[345]^x[344]^x[343]^x[340]^x[339]^x[338]^x[337]^x[334]^x[332]^x[329]^x[328]^x[327]^x[326]^x[324]^x[315]^x[314]^x[313]^x[304]^x[302]^x[248]^x[244]^x[233]^x[217]^x[211]^x[206]^x[200]^x[186]^x[185]^x[184]^x[183]^x[174]^x[172]^x[164]^x[142]^x[136]^x[130]^x[96]^x[90]^x[80]^x[78]^x[74]^x[73]^x[72]^x[69]^x[57]^x[46]^x[9]^x[7];
	y[13]=x[376]^x[365]^x[364]^x[353]^x[345]^x[344]^x[343]^x[342]^x[339]^x[338]^x[337]^x[336]^x[333]^x[331]^x[328]^x[327]^x[326]^x[325]^x[323]^x[314]^x[313]^x[312]^x[303]^x[301]^x[247]^x[243]^x[232]^x[216]^x[210]^x[205]^x[199]^x[185]^x[184]^x[183]^x[182]^x[173]^x[171]^x[163]^x[141]^x[135]^x[129]^x[89]^x[79]^x[77]^x[73]^x[72]^x[71]^x[68]^x[56]^x[45]^x[8]^x[6];
	y[12]=x[375]^x[364]^x[363]^x[352]^x[344]^x[343]^x[342]^x[338]^x[337]^x[336]^x[332]^x[327]^x[326]^x[325]^x[322]^x[313]^x[312]^x[311]^x[302]^x[300]^x[246]^x[242]^x[231]^x[215]^x[209]^x[204]^x[198]^x[184]^x[183]^x[182]^x[172]^x[162]^x[140]^x[134]^x[128]^x[88]^x[78]^x[76]^x[72]^x[71]^x[70]^x[67]^x[55]^x[44]^x[7]^x[5];
	y[11]=x[374]^x[363]^x[343]^x[342]^x[337]^x[336]^x[326]^x[325]^x[321]^x[320]^x[312]^x[311]^x[310]^x[301]^x[299]^x[246]^x[241]^x[235]^x[230]^x[214]^x[208]^x[203]^x[197]^x[183]^x[182]^x[161]^x[160]^x[139]^x[133]^x[87]^x[77]^x[75]^x[71]^x[70]^x[69]^x[66]^x[54]^x[43]^x[6]^x[5];
	y[10]=x[373]^x[362]^x[342]^x[341]^x[336]^x[335]^x[330]^x[325]^x[324]^x[320]^x[311]^x[310]^x[309]^x[300]^x[298]^x[240]^x[229]^x[213]^x[207]^x[202]^x[196]^x[182]^x[181]^x[170]^x[160]^x[138]^x[132]^x[86]^x[76]^x[74]^x[70]^x[69]^x[68]^x[65]^x[53]^x[42]^x[5];
	y[9]=x[372]^x[361]^x[351]^x[350]^x[345]^x[344]^x[341]^x[340]^x[339]^x[338]^x[335]^x[334]^x[333]^x[332]^x[330]^x[329]^x[327]^x[324]^x[323]^x[321]^x[310]^x[309]^x[308]^x[299]^x[297]^x[244]^x[243]^x[233]^x[212]^x[206]^x[201]^x[195]^x[191]^x[190]^x[181]^x[180]^x[179]^x[178]^x[170]^x[169]^x[167]^x[137]^x[131]^x[85]^x[79]^x[75]^x[73]^x[69]^x[67]^x[64]^x[52]^x[41];
	y[8]=x[371]^x[360]^x[350]^x[349]^x[344]^x[343]^x[340]^x[339]^x[338]^x[337]^x[334]^x[333]^x[332]^x[331]^x[329]^x[328]^x[326]^x[323]^x[322]^x[320]^x[309]^x[308]^x[307]^x[298]^x[296]^x[243]^x[242]^x[232]^x[211]^x[205]^x[200]^x[194]^x[190]^x[189]^x[180]^x[179]^x[178]^x[177]^x[169]^x[168]^x[166]^x[136]^x[130]^x[95]^x[89]^x[84]^x[78]^x[72]^x[66]^x[51]^x[40];
	y[7]=x[370]^x[359]^x[349]^x[348]^x[343]^x[342]^x[339]^x[338]^x[337]^x[336]^x[333]^x[332]^x[331]^x[328]^x[327]^x[325]^x[322]^x[321]^x[308]^x[307]^x[306]^x[297]^x[295]^x[242]^x[241]^x[231]^x[210]^x[204]^x[199]^x[193]^x[189]^x[188]^x[179]^x[178]^x[177]^x[176]^x[168]^x[167]^x[165]^x[135]^x[129]^x[94]^x[88]^x[83]^x[77]^x[71]^x[65]^x[50]^x[39];
	y[6]=x[369]^x[358]^x[348]^x[347]^x[342]^x[341]^x[338]^x[337]^x[336]^x[335]^x[332]^x[331]^x[330]^x[327]^x[326]^x[324]^x[321]^x[320]^x[307]^x[306]^x[305]^x[296]^x[294]^x[241]^x[240]^x[230]^x[209]^x[203]^x[198]^x[192]^x[188]^x[187]^x[178]^x[177]^x[176]^x[175]^x[167]^x[166]^x[164]^x[134]^x[128]^x[93]^x[87]^x[82]^x[76]^x[70]^x[64]^x[49]^x[38];
	y[5]=x[368]^x[357]^x[347]^x[346]^x[341]^x[340]^x[337]^x[336]^x[335]^x[334]^x[330]^x[329]^x[326]^x[325]^x[323]^x[306]^x[305]^x[304]^x[295]^x[293]^x[246]^x[239]^x[224]^x[208]^x[197]^x[187]^x[186]^x[177]^x[176]^x[175]^x[174]^x[166]^x[165]^x[163]^x[133]^x[92]^x[81]^x[75]^x[69]^x[64]^x[48]^x[37]^x[11]^x[0];
	y[4]=x[367]^x[356]^x[346]^x[345]^x[340]^x[339]^x[336]^x[335]^x[334]^x[333]^x[329]^x[328]^x[325]^x[324]^x[322]^x[305]^x[304]^x[303]^x[294]^x[292]^x[245]^x[238]^x[234]^x[207]^x[196]^x[186]^x[185]^x[176]^x[175]^x[174]^x[173]^x[165]^x[164]^x[162]^x[132]^x[91]^x[80]^x[68]^x[47]^x[36]^x[10];
	y[3]=x[366]^x[355]^x[345]^x[344]^x[339]^x[338]^x[335]^x[334]^x[333]^x[332]^x[328]^x[327]^x[324]^x[323]^x[321]^x[304]^x[303]^x[302]^x[293]^x[291]^x[244]^x[237]^x[233]^x[206]^x[195]^x[185]^x[184]^x[175]^x[174]^x[173]^x[172]^x[164]^x[163]^x[161]^x[131]^x[90]^x[79]^x[67]^x[46]^x[35]^x[9];
	y[2]=x[365]^x[354]^x[344]^x[343]^x[338]^x[337]^x[334]^x[333]^x[332]^x[331]^x[327]^x[326]^x[323]^x[322]^x[320]^x[303]^x[302]^x[301]^x[292]^x[290]^x[243]^x[236]^x[232]^x[205]^x[194]^x[184]^x[183]^x[174]^x[173]^x[172]^x[171]^x[163]^x[162]^x[160]^x[130]^x[89]^x[78]^x[66]^x[45]^x[34]^x[8];
	y[1]=x[364]^x[353]^x[343]^x[342]^x[337]^x[336]^x[333]^x[332]^x[331]^x[326]^x[325]^x[322]^x[321]^x[302]^x[301]^x[300]^x[291]^x[289]^x[242]^x[235]^x[231]^x[204]^x[193]^x[183]^x[182]^x[173]^x[172]^x[171]^x[162]^x[161]^x[129]^x[88]^x[77]^x[65]^x[44]^x[33]^x[7];
	y[0]=x[363]^x[352]^x[342]^x[336]^x[332]^x[331]^x[325]^x[321]^x[320]^x[301]^x[300]^x[299]^x[290]^x[288]^x[241]^x[235]^x[230]^x[224]^x[203]^x[192]^x[182]^x[172]^x[171]^x[161]^x[160]^x[128]^x[87]^x[76]^x[64]^x[43]^x[32]^x[6];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint51(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[378]^x[377]^x[368]^x[366]^x[357]^x[351]^x[350]^x[341]^x[339]^x[330]^x[317]^x[314]^x[311]^x[310]^x[308]^x[306]^x[304]^x[302]^x[300]^x[299]^x[298]^x[295]^x[293]^x[292]^x[289]^x[287]^x[279]^x[278]^x[277]^x[267]^x[266]^x[257]^x[223]^x[218]^x[213]^x[208]^x[202]^x[197]^x[191]^x[185]^x[181]^x[175]^x[170]^x[164]^x[157]^x[154]^x[150]^x[146]^x[142]^x[139]^x[138]^x[136]^x[135]^x[127]^x[121]^x[115]^x[109]^x[81]^x[63]^x[58]^x[57]^x[48]^x[44]^x[43]^x[38]^x[33]^x[31]^x[21]^x[10];
	y[30]=x[350]^x[349]^x[340]^x[338]^x[329]^x[318]^x[316]^x[312]^x[310]^x[309]^x[306]^x[305]^x[303]^x[300]^x[299]^x[298]^x[297]^x[295]^x[294]^x[292]^x[291]^x[289]^x[288]^x[286]^x[278]^x[277]^x[276]^x[266]^x[265]^x[256]^x[190]^x[184]^x[180]^x[174]^x[169]^x[163]^x[158]^x[156]^x[149]^x[146]^x[145]^x[138]^x[137]^x[135]^x[134]^x[126]^x[120]^x[114]^x[108]^x[80]^x[62]^x[56]^x[43]^x[42]^x[37]^x[36]^x[32]^x[30]^x[20]^x[9];
	y[29]=x[349]^x[348]^x[339]^x[337]^x[328]^x[317]^x[315]^x[311]^x[309]^x[308]^x[305]^x[304]^x[302]^x[298]^x[297]^x[296]^x[294]^x[293]^x[291]^x[290]^x[287]^x[285]^x[277]^x[276]^x[275]^x[266]^x[265]^x[264]^x[189]^x[183]^x[179]^x[173]^x[168]^x[162]^x[157]^x[155]^x[148]^x[145]^x[144]^x[137]^x[136]^x[134]^x[133]^x[125]^x[119]^x[113]^x[107]^x[79]^x[63]^x[61]^x[57]^x[55]^x[41]^x[35]^x[29]^x[19]^x[8];
	y[28]=x[348]^x[347]^x[338]^x[336]^x[327]^x[316]^x[314]^x[310]^x[308]^x[307]^x[304]^x[303]^x[301]^x[297]^x[296]^x[295]^x[293]^x[292]^x[290]^x[289]^x[286]^x[284]^x[276]^x[275]^x[274]^x[265]^x[264]^x[263]^x[188]^x[182]^x[178]^x[172]^x[167]^x[161]^x[156]^x[154]^x[147]^x[144]^x[143]^x[136]^x[135]^x[133]^x[132]^x[124]^x[118]^x[112]^x[106]^x[78]^x[62]^x[60]^x[56]^x[54]^x[40]^x[34]^x[28]^x[18]^x[7];
	y[27]=x[347]^x[346]^x[337]^x[335]^x[326]^x[315]^x[313]^x[309]^x[307]^x[306]^x[303]^x[302]^x[300]^x[296]^x[295]^x[294]^x[292]^x[291]^x[289]^x[288]^x[285]^x[283]^x[275]^x[274]^x[273]^x[264]^x[263]^x[262]^x[187]^x[181]^x[177]^x[171]^x[166]^x[160]^x[155]^x[153]^x[146]^x[143]^x[142]^x[135]^x[134]^x[132]^x[131]^x[123]^x[117]^x[111]^x[105]^x[77]^x[61]^x[59]^x[55]^x[53]^x[39]^x[33]^x[27]^x[17]^x[6];
	y[26]=x[383]^x[382]^x[373]^x[372]^x[371]^x[363]^x[352]^x[346]^x[345]^x[336]^x[334]^x[325]^x[317]^x[314]^x[312]^x[309]^x[307]^x[306]^x[305]^x[302]^x[301]^x[299]^x[297]^x[294]^x[293]^x[291]^x[290]^x[288]^x[284]^x[282]^x[274]^x[273]^x[272]^x[263]^x[262]^x[261]^x[218]^x[213]^x[207]^x[203]^x[192]^x[191]^x[186]^x[180]^x[176]^x[165]^x[154]^x[152]^x[149]^x[148]^x[147]^x[145]^x[143]^x[134]^x[133]^x[131]^x[130]^x[122]^x[116]^x[110]^x[104]^x[76]^x[60]^x[58]^x[54]^x[53]^x[52]^x[43]^x[38]^x[26]^x[16]^x[5];
	y[25]=x[381]^x[372]^x[370]^x[345]^x[344]^x[335]^x[333]^x[324]^x[319]^x[316]^x[313]^x[311]^x[308]^x[306]^x[305]^x[304]^x[301]^x[300]^x[296]^x[293]^x[292]^x[290]^x[289]^x[283]^x[281]^x[273]^x[272]^x[271]^x[262]^x[261]^x[260]^x[212]^x[206]^x[190]^x[185]^x[179]^x[175]^x[164]^x[159]^x[151]^x[148]^x[146]^x[144]^x[142]^x[141]^x[138]^x[133]^x[130]^x[129]^x[121]^x[115]^x[109]^x[103]^x[75]^x[59]^x[57]^x[53]^x[52]^x[51]^x[37]^x[25]^x[15]^x[4];
	y[24]=x[380]^x[371]^x[369]^x[344]^x[343]^x[334]^x[332]^x[323]^x[318]^x[315]^x[312]^x[310]^x[307]^x[305]^x[304]^x[303]^x[300]^x[299]^x[295]^x[292]^x[291]^x[289]^x[288]^x[282]^x[280]^x[272]^x[271]^x[270]^x[261]^x[260]^x[259]^x[211]^x[205]^x[189]^x[184]^x[178]^x[174]^x[163]^x[158]^x[150]^x[147]^x[145]^x[143]^x[141]^x[140]^x[137]^x[132]^x[129]^x[128]^x[120]^x[114]^x[108]^x[102]^x[74]^x[58]^x[56]^x[52]^x[51]^x[50]^x[36]^x[24]^x[14]^x[3];
	y[23]=x[379]^x[370]^x[368]^x[343]^x[342]^x[333]^x[331]^x[322]^x[317]^x[314]^x[311]^x[306]^x[304]^x[302]^x[294]^x[292]^x[291]^x[290]^x[281]^x[279]^x[271]^x[270]^x[269]^x[260]^x[259]^x[258]^x[210]^x[204]^x[188]^x[183]^x[177]^x[173]^x[162]^x[157]^x[146]^x[144]^x[142]^x[140]^x[138]^x[136]^x[131]^x[119]^x[113]^x[107]^x[101]^x[73]^x[57]^x[55]^x[51]^x[50]^x[49]^x[35]^x[23]^x[13]^x[2];
	y[22]=x[378]^x[369]^x[367]^x[342]^x[341]^x[332]^x[330]^x[321]^x[316]^x[313]^x[310]^x[305]^x[303]^x[301]^x[293]^x[291]^x[290]^x[289]^x[280]^x[278]^x[270]^x[269]^x[268]^x[259]^x[258]^x[257]^x[209]^x[203]^x[187]^x[182]^x[176]^x[172]^x[161]^x[156]^x[145]^x[143]^x[141]^x[139]^x[137]^x[135]^x[130]^x[118]^x[112]^x[106]^x[100]^x[72]^x[56]^x[54]^x[50]^x[49]^x[48]^x[34]^x[22]^x[12]^x[1];
	y[21]=x[377]^x[368]^x[366]^x[341]^x[340]^x[331]^x[329]^x[320]^x[315]^x[312]^x[304]^x[303]^x[302]^x[300]^x[298]^x[290]^x[289]^x[288]^x[279]^x[277]^x[269]^x[268]^x[267]^x[258]^x[257]^x[256]^x[208]^x[203]^x[192]^x[186]^x[181]^x[175]^x[171]^x[160]^x[155]^x[149]^x[144]^x[142]^x[140]^x[136]^x[134]^x[129]^x[117]^x[111]^x[105]^x[99]^x[71]^x[55]^x[53]^x[49]^x[48]^x[47]^x[33]^x[21]^x[11]^x[0];
	y[20]=x[378]^x[377]^x[366]^x[351]^x[340]^x[339]^x[328]^x[319]^x[318]^x[317]^x[314]^x[313]^x[312]^x[311]^x[308]^x[306]^x[302]^x[300]^x[299]^x[298]^x[292]^x[288]^x[287]^x[278]^x[276]^x[268]^x[267]^x[257]^x[256]^x[223]^x[222]^x[218]^x[201]^x[191]^x[185]^x[180]^x[174]^x[159]^x[158]^x[157]^x[154]^x[146]^x[142]^x[139]^x[138]^x[136]^x[133]^x[128]^x[116]^x[110]^x[104]^x[98]^x[70]^x[58]^x[54]^x[52]^x[48]^x[46]^x[32]^x[31]^x[20];
	y[19]=x[350]^x[339]^x[338]^x[327]^x[319]^x[318]^x[317]^x[316]^x[313]^x[312]^x[311]^x[310]^x[307]^x[305]^x[301]^x[299]^x[297]^x[291]^x[287]^x[286]^x[277]^x[275]^x[267]^x[256]^x[221]^x[211]^x[200]^x[190]^x[184]^x[179]^x[173]^x[159]^x[158]^x[157]^x[156]^x[147]^x[145]^x[137]^x[115]^x[109]^x[103]^x[97]^x[69]^x[63]^x[57]^x[53]^x[51]^x[47]^x[45]^x[42]^x[36]^x[30]^x[19];
	y[18]=x[349]^x[338]^x[337]^x[326]^x[318]^x[317]^x[316]^x[315]^x[312]^x[311]^x[310]^x[309]^x[306]^x[304]^x[300]^x[298]^x[296]^x[290]^x[287]^x[286]^x[285]^x[276]^x[274]^x[220]^x[210]^x[199]^x[189]^x[183]^x[178]^x[172]^x[158]^x[157]^x[156]^x[155]^x[146]^x[144]^x[136]^x[114]^x[108]^x[102]^x[96]^x[68]^x[62]^x[56]^x[52]^x[50]^x[46]^x[44]^x[41]^x[35]^x[29]^x[18];
	y[17]=x[374]^x[373]^x[362]^x[352]^x[348]^x[337]^x[336]^x[325]^x[317]^x[316]^x[315]^x[314]^x[311]^x[310]^x[309]^x[308]^x[305]^x[303]^x[298]^x[297]^x[295]^x[289]^x[288]^x[286]^x[285]^x[284]^x[275]^x[273]^x[219]^x[209]^x[198]^x[188]^x[182]^x[177]^x[171]^x[157]^x[156]^x[155]^x[154]^x[145]^x[143]^x[139]^x[138]^x[135]^x[133]^x[132]^x[128]^x[113]^x[107]^x[101]^x[67]^x[61]^x[55]^x[51]^x[49]^x[45]^x[43]^x[40]^x[34]^x[28]^x[17];
	y[16]=x[372]^x[361]^x[347]^x[336]^x[335]^x[324]^x[316]^x[315]^x[314]^x[313]^x[310]^x[309]^x[308]^x[307]^x[304]^x[302]^x[298]^x[297]^x[296]^x[294]^x[288]^x[285]^x[284]^x[283]^x[274]^x[272]^x[218]^x[208]^x[197]^x[187]^x[181]^x[176]^x[170]^x[156]^x[155]^x[154]^x[153]^x[144]^x[142]^x[137]^x[134]^x[131]^x[112]^x[106]^x[100]^x[66]^x[60]^x[54]^x[50]^x[48]^x[44]^x[42]^x[39]^x[33]^x[27]^x[16];
	y[15]=x[373]^x[371]^x[362]^x[360]^x[346]^x[335]^x[334]^x[323]^x[315]^x[314]^x[313]^x[312]^x[309]^x[308]^x[307]^x[306]^x[303]^x[301]^x[298]^x[297]^x[296]^x[295]^x[293]^x[284]^x[283]^x[282]^x[273]^x[271]^x[217]^x[213]^x[202]^x[186]^x[180]^x[175]^x[169]^x[155]^x[154]^x[153]^x[152]^x[143]^x[141]^x[138]^x[136]^x[133]^x[132]^x[130]^x[111]^x[105]^x[99]^x[65]^x[59]^x[49]^x[47]^x[43]^x[42]^x[41]^x[38]^x[32]^x[26]^x[15];
	y[14]=x[372]^x[370]^x[361]^x[359]^x[345]^x[334]^x[333]^x[322]^x[314]^x[313]^x[312]^x[311]^x[308]^x[307]^x[306]^x[305]^x[302]^x[300]^x[297]^x[296]^x[295]^x[294]^x[292]^x[283]^x[282]^x[281]^x[272]^x[270]^x[216]^x[212]^x[201]^x[185]^x[179]^x[174]^x[168]^x[154]^x[153]^x[152]^x[151]^x[142]^x[140]^x[137]^x[135]^x[132]^x[131]^x[129]^x[110]^x[104]^x[98]^x[64]^x[58]^x[48]^x[46]^x[42]^x[41]^x[40]^x[37]^x[25]^x[14];
	y[13]=x[371]^x[369]^x[360]^x[358]^x[344]^x[333]^x[332]^x[321]^x[313]^x[312]^x[311]^x[310]^x[307]^x[306]^x[305]^x[304]^x[301]^x[299]^x[296]^x[295]^x[294]^x[293]^x[291]^x[282]^x[281]^x[280]^x[271]^x[269]^x[215]^x[211]^x[200]^x[184]^x[178]^x[173]^x[167]^x[153]^x[152]^x[151]^x[150]^x[141]^x[139]^x[136]^x[134]^x[131]^x[130]^x[128]^x[109]^x[103]^x[97]^x[57]^x[47]^x[45]^x[41]^x[40]^x[39]^x[36]^x[24]^x[13];
	y[12]=x[370]^x[368]^x[359]^x[357]^x[343]^x[332]^x[331]^x[320]^x[312]^x[311]^x[310]^x[306]^x[305]^x[304]^x[300]^x[295]^x[294]^x[293]^x[290]^x[281]^x[280]^x[279]^x[270]^x[268]^x[214]^x[210]^x[199]^x[183]^x[177]^x[172]^x[166]^x[152]^x[151]^x[150]^x[140]^x[135]^x[133]^x[130]^x[129]^x[108]^x[102]^x[96]^x[56]^x[46]^x[44]^x[40]^x[39]^x[38]^x[35]^x[23]^x[12];
	y[11]=x[369]^x[368]^x[358]^x[357]^x[342]^x[331]^x[311]^x[310]^x[305]^x[304]^x[294]^x[293]^x[289]^x[288]^x[280]^x[279]^x[278]^x[269]^x[267]^x[214]^x[209]^x[203]^x[198]^x[182]^x[176]^x[171]^x[165]^x[151]^x[150]^x[134]^x[133]^x[129]^x[107]^x[101]^x[55]^x[45]^x[43]^x[39]^x[38]^x[37]^x[34]^x[22]^x[11];
	y[10]=x[368]^x[357]^x[341]^x[330]^x[310]^x[309]^x[304]^x[303]^x[298]^x[293]^x[292]^x[288]^x[279]^x[278]^x[277]^x[268]^x[266]^x[208]^x[197]^x[181]^x[175]^x[170]^x[164]^x[150]^x[149]^x[138]^x[133]^x[128]^x[106]^x[100]^x[54]^x[44]^x[42]^x[38]^x[37]^x[36]^x[33]^x[21]^x[10];
	y[9]=x[340]^x[329]^x[319]^x[318]^x[313]^x[312]^x[309]^x[308]^x[307]^x[306]^x[303]^x[302]^x[301]^x[300]^x[298]^x[297]^x[295]^x[292]^x[291]^x[289]^x[278]^x[277]^x[276]^x[267]^x[265]^x[212]^x[211]^x[201]^x[180]^x[174]^x[169]^x[163]^x[159]^x[158]^x[149]^x[148]^x[147]^x[146]^x[138]^x[137]^x[135]^x[105]^x[99]^x[53]^x[47]^x[43]^x[41]^x[37]^x[35]^x[32]^x[20]^x[9];
	y[8]=x[339]^x[328]^x[318]^x[317]^x[312]^x[311]^x[308]^x[307]^x[306]^x[305]^x[302]^x[301]^x[300]^x[299]^x[297]^x[296]^x[294]^x[291]^x[290]^x[288]^x[277]^x[276]^x[275]^x[266]^x[264]^x[211]^x[210]^x[200]^x[179]^x[173]^x[168]^x[162]^x[158]^x[157]^x[148]^x[147]^x[146]^x[145]^x[137]^x[136]^x[134]^x[104]^x[98]^x[63]^x[57]^x[52]^x[46]^x[40]^x[34]^x[19]^x[8];
	y[7]=x[338]^x[327]^x[317]^x[316]^x[311]^x[310]^x[307]^x[306]^x[305]^x[304]^x[301]^x[300]^x[299]^x[296]^x[295]^x[293]^x[290]^x[289]^x[276]^x[275]^x[274]^x[265]^x[263]^x[210]^x[209]^x[199]^x[178]^x[172]^x[167]^x[161]^x[157]^x[156]^x[147]^x[146]^x[145]^x[144]^x[136]^x[135]^x[133]^x[103]^x[97]^x[62]^x[56]^x[51]^x[45]^x[39]^x[33]^x[18]^x[7];
	y[6]=x[337]^x[326]^x[316]^x[315]^x[310]^x[309]^x[306]^x[305]^x[304]^x[303]^x[300]^x[299]^x[298]^x[295]^x[294]^x[292]^x[289]^x[288]^x[275]^x[274]^x[273]^x[264]^x[262]^x[209]^x[208]^x[198]^x[177]^x[171]^x[166]^x[160]^x[156]^x[155]^x[146]^x[145]^x[144]^x[143]^x[135]^x[134]^x[132]^x[102]^x[96]^x[61]^x[55]^x[50]^x[44]^x[38]^x[32]^x[17]^x[6];
	y[5]=x[374]^x[352]^x[336]^x[325]^x[315]^x[314]^x[309]^x[308]^x[305]^x[304]^x[303]^x[302]^x[298]^x[297]^x[294]^x[293]^x[291]^x[274]^x[273]^x[272]^x[263]^x[261]^x[214]^x[207]^x[192]^x[176]^x[165]^x[155]^x[154]^x[145]^x[144]^x[143]^x[142]^x[139]^x[134]^x[131]^x[128]^x[101]^x[60]^x[49]^x[43]^x[37]^x[32]^x[16]^x[5];
	y[4]=x[373]^x[362]^x[335]^x[324]^x[314]^x[313]^x[308]^x[307]^x[304]^x[303]^x[302]^x[301]^x[297]^x[296]^x[293]^x[292]^x[290]^x[273]^x[272]^x[271]^x[262]^x[260]^x[213]^x[206]^x[202]^x[175]^x[164]^x[154]^x[153]^x[144]^x[143]^x[142]^x[141]^x[138]^x[133]^x[130]^x[100]^x[59]^x[48]^x[36]^x[15]^x[4];
	y[3]=x[372]^x[361]^x[334]^x[323]^x[313]^x[312]^x[307]^x[306]^x[303]^x[302]^x[301]^x[300]^x[296]^x[295]^x[292]^x[291]^x[289]^x[272]^x[271]^x[270]^x[261]^x[259]^x[212]^x[205]^x[201]^x[174]^x[163]^x[153]^x[152]^x[143]^x[142]^x[141]^x[140]^x[137]^x[132]^x[129]^x[99]^x[58]^x[47]^x[35]^x[14]^x[3];
	y[2]=x[371]^x[360]^x[333]^x[322]^x[312]^x[311]^x[306]^x[305]^x[302]^x[301]^x[300]^x[299]^x[295]^x[294]^x[291]^x[290]^x[288]^x[271]^x[270]^x[269]^x[260]^x[258]^x[211]^x[204]^x[200]^x[173]^x[162]^x[152]^x[151]^x[142]^x[141]^x[140]^x[139]^x[136]^x[131]^x[128]^x[98]^x[57]^x[46]^x[34]^x[13]^x[2];
	y[1]=x[370]^x[359]^x[332]^x[321]^x[311]^x[310]^x[305]^x[304]^x[301]^x[300]^x[299]^x[294]^x[293]^x[290]^x[289]^x[270]^x[269]^x[268]^x[259]^x[257]^x[210]^x[203]^x[199]^x[172]^x[161]^x[151]^x[150]^x[141]^x[140]^x[139]^x[135]^x[130]^x[97]^x[56]^x[45]^x[33]^x[12]^x[1];
	y[0]=x[369]^x[358]^x[331]^x[320]^x[310]^x[304]^x[300]^x[299]^x[293]^x[289]^x[288]^x[269]^x[268]^x[267]^x[258]^x[256]^x[209]^x[203]^x[198]^x[192]^x[171]^x[160]^x[150]^x[140]^x[139]^x[134]^x[129]^x[96]^x[55]^x[44]^x[32]^x[11]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint52(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[373]^x[363]^x[352]^x[346]^x[345]^x[336]^x[334]^x[325]^x[319]^x[318]^x[309]^x[307]^x[298]^x[285]^x[282]^x[279]^x[278]^x[276]^x[274]^x[272]^x[270]^x[268]^x[267]^x[266]^x[263]^x[261]^x[260]^x[257]^x[255]^x[247]^x[246]^x[245]^x[235]^x[234]^x[225]^x[191]^x[186]^x[181]^x[176]^x[170]^x[165]^x[125]^x[122]^x[118]^x[114]^x[110]^x[107]^x[106]^x[104]^x[103]^x[95]^x[89]^x[83]^x[77]^x[49]^x[31]^x[26]^x[25]^x[16]^x[12]^x[11]^x[6]^x[1];
	y[30]=x[383]^x[382]^x[372]^x[318]^x[317]^x[308]^x[306]^x[297]^x[286]^x[284]^x[280]^x[278]^x[277]^x[274]^x[273]^x[271]^x[268]^x[267]^x[266]^x[265]^x[263]^x[262]^x[260]^x[259]^x[257]^x[256]^x[254]^x[246]^x[245]^x[244]^x[234]^x[233]^x[224]^x[126]^x[124]^x[117]^x[114]^x[113]^x[106]^x[105]^x[103]^x[102]^x[94]^x[88]^x[82]^x[76]^x[48]^x[30]^x[24]^x[11]^x[10]^x[5]^x[4]^x[0];
	y[29]=x[382]^x[381]^x[371]^x[317]^x[316]^x[307]^x[305]^x[296]^x[285]^x[283]^x[279]^x[277]^x[276]^x[273]^x[272]^x[270]^x[266]^x[265]^x[264]^x[262]^x[261]^x[259]^x[258]^x[255]^x[253]^x[245]^x[244]^x[243]^x[234]^x[233]^x[232]^x[125]^x[123]^x[116]^x[113]^x[112]^x[105]^x[104]^x[102]^x[101]^x[93]^x[87]^x[81]^x[75]^x[47]^x[31]^x[29]^x[25]^x[23]^x[9]^x[3];
	y[28]=x[381]^x[380]^x[370]^x[316]^x[315]^x[306]^x[304]^x[295]^x[284]^x[282]^x[278]^x[276]^x[275]^x[272]^x[271]^x[269]^x[265]^x[264]^x[263]^x[261]^x[260]^x[258]^x[257]^x[254]^x[252]^x[244]^x[243]^x[242]^x[233]^x[232]^x[231]^x[124]^x[122]^x[115]^x[112]^x[111]^x[104]^x[103]^x[101]^x[100]^x[92]^x[86]^x[80]^x[74]^x[46]^x[30]^x[28]^x[24]^x[22]^x[8]^x[2];
	y[27]=x[380]^x[379]^x[369]^x[315]^x[314]^x[305]^x[303]^x[294]^x[283]^x[281]^x[277]^x[275]^x[274]^x[271]^x[270]^x[268]^x[264]^x[263]^x[262]^x[260]^x[259]^x[257]^x[256]^x[253]^x[251]^x[243]^x[242]^x[241]^x[232]^x[231]^x[230]^x[123]^x[121]^x[114]^x[111]^x[110]^x[103]^x[102]^x[100]^x[99]^x[91]^x[85]^x[79]^x[73]^x[45]^x[29]^x[27]^x[23]^x[21]^x[7]^x[1];
	y[26]=x[379]^x[378]^x[368]^x[351]^x[350]^x[341]^x[340]^x[339]^x[331]^x[320]^x[314]^x[313]^x[304]^x[302]^x[293]^x[285]^x[282]^x[280]^x[277]^x[275]^x[274]^x[273]^x[270]^x[269]^x[267]^x[265]^x[262]^x[261]^x[259]^x[258]^x[256]^x[252]^x[250]^x[242]^x[241]^x[240]^x[231]^x[230]^x[229]^x[186]^x[181]^x[175]^x[171]^x[160]^x[159]^x[138]^x[122]^x[120]^x[117]^x[116]^x[115]^x[113]^x[111]^x[102]^x[101]^x[99]^x[98]^x[90]^x[84]^x[78]^x[72]^x[44]^x[28]^x[26]^x[22]^x[21]^x[20]^x[11]^x[6];
	y[25]=x[378]^x[377]^x[367]^x[349]^x[340]^x[338]^x[313]^x[312]^x[303]^x[301]^x[292]^x[287]^x[284]^x[281]^x[279]^x[276]^x[274]^x[273]^x[272]^x[269]^x[268]^x[264]^x[261]^x[260]^x[258]^x[257]^x[251]^x[249]^x[241]^x[240]^x[239]^x[230]^x[229]^x[228]^x[180]^x[174]^x[158]^x[137]^x[127]^x[119]^x[116]^x[114]^x[112]^x[110]^x[109]^x[106]^x[101]^x[98]^x[97]^x[89]^x[83]^x[77]^x[71]^x[43]^x[27]^x[25]^x[21]^x[20]^x[19]^x[5];
	y[24]=x[377]^x[376]^x[366]^x[348]^x[339]^x[337]^x[312]^x[311]^x[302]^x[300]^x[291]^x[286]^x[283]^x[280]^x[278]^x[275]^x[273]^x[272]^x[271]^x[268]^x[267]^x[263]^x[260]^x[259]^x[257]^x[256]^x[250]^x[248]^x[240]^x[239]^x[238]^x[229]^x[228]^x[227]^x[179]^x[173]^x[157]^x[136]^x[126]^x[118]^x[115]^x[113]^x[111]^x[109]^x[108]^x[105]^x[100]^x[97]^x[96]^x[88]^x[82]^x[76]^x[70]^x[42]^x[26]^x[24]^x[20]^x[19]^x[18]^x[4];
	y[23]=x[376]^x[375]^x[365]^x[347]^x[338]^x[336]^x[311]^x[310]^x[301]^x[299]^x[290]^x[285]^x[282]^x[279]^x[274]^x[272]^x[270]^x[262]^x[260]^x[259]^x[258]^x[249]^x[247]^x[239]^x[238]^x[237]^x[228]^x[227]^x[226]^x[178]^x[172]^x[156]^x[135]^x[125]^x[114]^x[112]^x[110]^x[108]^x[106]^x[104]^x[99]^x[87]^x[81]^x[75]^x[69]^x[41]^x[25]^x[23]^x[19]^x[18]^x[17]^x[3];
	y[22]=x[375]^x[374]^x[364]^x[346]^x[337]^x[335]^x[310]^x[309]^x[300]^x[298]^x[289]^x[284]^x[281]^x[278]^x[273]^x[271]^x[269]^x[261]^x[259]^x[258]^x[257]^x[248]^x[246]^x[238]^x[237]^x[236]^x[227]^x[226]^x[225]^x[177]^x[171]^x[155]^x[134]^x[124]^x[113]^x[111]^x[109]^x[107]^x[105]^x[103]^x[98]^x[86]^x[80]^x[74]^x[68]^x[40]^x[24]^x[22]^x[18]^x[17]^x[16]^x[2];
	y[21]=x[374]^x[373]^x[363]^x[345]^x[336]^x[334]^x[309]^x[308]^x[299]^x[297]^x[288]^x[283]^x[280]^x[272]^x[271]^x[270]^x[268]^x[266]^x[258]^x[257]^x[256]^x[247]^x[245]^x[237]^x[236]^x[235]^x[226]^x[225]^x[224]^x[176]^x[171]^x[160]^x[154]^x[133]^x[123]^x[117]^x[112]^x[110]^x[108]^x[104]^x[102]^x[97]^x[85]^x[79]^x[73]^x[67]^x[39]^x[23]^x[21]^x[17]^x[16]^x[15]^x[1];
	y[20]=x[373]^x[372]^x[362]^x[346]^x[345]^x[334]^x[319]^x[308]^x[307]^x[296]^x[287]^x[286]^x[285]^x[282]^x[281]^x[280]^x[279]^x[276]^x[274]^x[270]^x[268]^x[267]^x[266]^x[260]^x[256]^x[255]^x[246]^x[244]^x[236]^x[235]^x[225]^x[224]^x[191]^x[190]^x[186]^x[169]^x[127]^x[126]^x[125]^x[122]^x[114]^x[110]^x[107]^x[106]^x[104]^x[101]^x[96]^x[84]^x[78]^x[72]^x[66]^x[38]^x[26]^x[22]^x[20]^x[16]^x[14]^x[0];
	y[19]=x[372]^x[371]^x[361]^x[318]^x[307]^x[306]^x[295]^x[287]^x[286]^x[285]^x[284]^x[281]^x[280]^x[279]^x[278]^x[275]^x[273]^x[269]^x[267]^x[265]^x[259]^x[255]^x[254]^x[245]^x[243]^x[235]^x[224]^x[189]^x[179]^x[168]^x[127]^x[126]^x[125]^x[124]^x[115]^x[113]^x[105]^x[83]^x[77]^x[71]^x[65]^x[37]^x[31]^x[25]^x[21]^x[19]^x[15]^x[13]^x[10]^x[4];
	y[18]=x[371]^x[370]^x[360]^x[317]^x[306]^x[305]^x[294]^x[286]^x[285]^x[284]^x[283]^x[280]^x[279]^x[278]^x[277]^x[274]^x[272]^x[268]^x[266]^x[264]^x[258]^x[255]^x[254]^x[253]^x[244]^x[242]^x[188]^x[178]^x[167]^x[126]^x[125]^x[124]^x[123]^x[114]^x[112]^x[104]^x[82]^x[76]^x[70]^x[64]^x[36]^x[30]^x[24]^x[20]^x[18]^x[14]^x[12]^x[9]^x[3];
	y[17]=x[370]^x[369]^x[359]^x[342]^x[341]^x[330]^x[320]^x[316]^x[305]^x[304]^x[293]^x[285]^x[284]^x[283]^x[282]^x[279]^x[278]^x[277]^x[276]^x[273]^x[271]^x[266]^x[265]^x[263]^x[257]^x[256]^x[254]^x[253]^x[252]^x[243]^x[241]^x[187]^x[177]^x[166]^x[125]^x[124]^x[123]^x[122]^x[113]^x[111]^x[107]^x[106]^x[103]^x[101]^x[100]^x[96]^x[81]^x[75]^x[69]^x[35]^x[29]^x[23]^x[19]^x[17]^x[13]^x[11]^x[8]^x[2];
	y[16]=x[369]^x[368]^x[358]^x[340]^x[329]^x[315]^x[304]^x[303]^x[292]^x[284]^x[283]^x[282]^x[281]^x[278]^x[277]^x[276]^x[275]^x[272]^x[270]^x[266]^x[265]^x[264]^x[262]^x[256]^x[253]^x[252]^x[251]^x[242]^x[240]^x[186]^x[176]^x[165]^x[124]^x[123]^x[122]^x[121]^x[112]^x[110]^x[105]^x[102]^x[99]^x[80]^x[74]^x[68]^x[34]^x[28]^x[22]^x[18]^x[16]^x[12]^x[10]^x[7]^x[1];
	y[15]=x[368]^x[367]^x[357]^x[341]^x[339]^x[330]^x[328]^x[314]^x[303]^x[302]^x[291]^x[283]^x[282]^x[281]^x[280]^x[277]^x[276]^x[275]^x[274]^x[271]^x[269]^x[266]^x[265]^x[264]^x[263]^x[261]^x[252]^x[251]^x[250]^x[241]^x[239]^x[185]^x[181]^x[170]^x[123]^x[122]^x[121]^x[120]^x[111]^x[109]^x[106]^x[104]^x[101]^x[100]^x[98]^x[79]^x[73]^x[67]^x[33]^x[27]^x[17]^x[15]^x[11]^x[10]^x[9]^x[6]^x[0];
	y[14]=x[367]^x[366]^x[356]^x[340]^x[338]^x[329]^x[327]^x[313]^x[302]^x[301]^x[290]^x[282]^x[281]^x[280]^x[279]^x[276]^x[275]^x[274]^x[273]^x[270]^x[268]^x[265]^x[264]^x[263]^x[262]^x[260]^x[251]^x[250]^x[249]^x[240]^x[238]^x[184]^x[180]^x[169]^x[122]^x[121]^x[120]^x[119]^x[110]^x[108]^x[105]^x[103]^x[100]^x[99]^x[97]^x[78]^x[72]^x[66]^x[32]^x[26]^x[16]^x[14]^x[10]^x[9]^x[8]^x[5];
	y[13]=x[366]^x[365]^x[355]^x[339]^x[337]^x[328]^x[326]^x[312]^x[301]^x[300]^x[289]^x[281]^x[280]^x[279]^x[278]^x[275]^x[274]^x[273]^x[272]^x[269]^x[267]^x[264]^x[263]^x[262]^x[261]^x[259]^x[250]^x[249]^x[248]^x[239]^x[237]^x[183]^x[179]^x[168]^x[121]^x[120]^x[119]^x[118]^x[109]^x[107]^x[104]^x[102]^x[99]^x[98]^x[96]^x[77]^x[71]^x[65]^x[25]^x[15]^x[13]^x[9]^x[8]^x[7]^x[4];
	y[12]=x[365]^x[364]^x[354]^x[338]^x[336]^x[327]^x[325]^x[311]^x[300]^x[299]^x[288]^x[280]^x[279]^x[278]^x[274]^x[273]^x[272]^x[268]^x[263]^x[262]^x[261]^x[258]^x[249]^x[248]^x[247]^x[238]^x[236]^x[182]^x[178]^x[167]^x[120]^x[119]^x[118]^x[108]^x[103]^x[101]^x[98]^x[97]^x[76]^x[70]^x[64]^x[24]^x[14]^x[12]^x[8]^x[7]^x[6]^x[3];
	y[11]=x[364]^x[363]^x[353]^x[337]^x[336]^x[326]^x[325]^x[310]^x[299]^x[279]^x[278]^x[273]^x[272]^x[262]^x[261]^x[257]^x[256]^x[248]^x[247]^x[246]^x[237]^x[235]^x[182]^x[177]^x[171]^x[166]^x[119]^x[118]^x[102]^x[101]^x[97]^x[75]^x[69]^x[23]^x[13]^x[11]^x[7]^x[6]^x[5]^x[2];
	y[10]=x[363]^x[362]^x[352]^x[336]^x[325]^x[309]^x[298]^x[278]^x[277]^x[272]^x[271]^x[266]^x[261]^x[260]^x[256]^x[247]^x[246]^x[245]^x[236]^x[234]^x[176]^x[165]^x[118]^x[117]^x[106]^x[101]^x[96]^x[74]^x[68]^x[22]^x[12]^x[10]^x[6]^x[5]^x[4]^x[1];
	y[9]=x[383]^x[361]^x[308]^x[297]^x[287]^x[286]^x[281]^x[280]^x[277]^x[276]^x[275]^x[274]^x[271]^x[270]^x[269]^x[268]^x[266]^x[265]^x[263]^x[260]^x[259]^x[257]^x[246]^x[245]^x[244]^x[235]^x[233]^x[180]^x[179]^x[169]^x[127]^x[126]^x[117]^x[116]^x[115]^x[114]^x[106]^x[105]^x[103]^x[73]^x[67]^x[21]^x[15]^x[11]^x[9]^x[5]^x[3]^x[0];
	y[8]=x[382]^x[360]^x[307]^x[296]^x[286]^x[285]^x[280]^x[279]^x[276]^x[275]^x[274]^x[273]^x[270]^x[269]^x[268]^x[267]^x[265]^x[264]^x[262]^x[259]^x[258]^x[256]^x[245]^x[244]^x[243]^x[234]^x[232]^x[179]^x[178]^x[168]^x[126]^x[125]^x[116]^x[115]^x[114]^x[113]^x[105]^x[104]^x[102]^x[72]^x[66]^x[31]^x[25]^x[20]^x[14]^x[8]^x[2];
	y[7]=x[381]^x[359]^x[306]^x[295]^x[285]^x[284]^x[279]^x[278]^x[275]^x[274]^x[273]^x[272]^x[269]^x[268]^x[267]^x[264]^x[263]^x[261]^x[258]^x[257]^x[244]^x[243]^x[242]^x[233]^x[231]^x[178]^x[177]^x[167]^x[125]^x[124]^x[115]^x[114]^x[113]^x[112]^x[104]^x[103]^x[101]^x[71]^x[65]^x[30]^x[24]^x[19]^x[13]^x[7]^x[1];
	y[6]=x[380]^x[358]^x[305]^x[294]^x[284]^x[283]^x[278]^x[277]^x[274]^x[273]^x[272]^x[271]^x[268]^x[267]^x[266]^x[263]^x[262]^x[260]^x[257]^x[256]^x[243]^x[242]^x[241]^x[232]^x[230]^x[177]^x[176]^x[166]^x[124]^x[123]^x[114]^x[113]^x[112]^x[111]^x[103]^x[102]^x[100]^x[70]^x[64]^x[29]^x[23]^x[18]^x[12]^x[6]^x[0];
	y[5]=x[379]^x[357]^x[342]^x[320]^x[304]^x[293]^x[283]^x[282]^x[277]^x[276]^x[273]^x[272]^x[271]^x[270]^x[266]^x[265]^x[262]^x[261]^x[259]^x[242]^x[241]^x[240]^x[231]^x[229]^x[182]^x[175]^x[160]^x[138]^x[123]^x[122]^x[113]^x[112]^x[111]^x[110]^x[107]^x[102]^x[99]^x[96]^x[69]^x[28]^x[17]^x[11]^x[5]^x[0];
	y[4]=x[378]^x[356]^x[341]^x[330]^x[303]^x[292]^x[282]^x[281]^x[276]^x[275]^x[272]^x[271]^x[270]^x[269]^x[265]^x[264]^x[261]^x[260]^x[258]^x[241]^x[240]^x[239]^x[230]^x[228]^x[181]^x[174]^x[170]^x[137]^x[122]^x[121]^x[112]^x[111]^x[110]^x[109]^x[106]^x[101]^x[98]^x[68]^x[27]^x[16]^x[4];
	y[3]=x[377]^x[355]^x[340]^x[329]^x[302]^x[291]^x[281]^x[280]^x[275]^x[274]^x[271]^x[270]^x[269]^x[268]^x[264]^x[263]^x[260]^x[259]^x[257]^x[240]^x[239]^x[238]^x[229]^x[227]^x[180]^x[173]^x[169]^x[136]^x[121]^x[120]^x[111]^x[110]^x[109]^x[108]^x[105]^x[100]^x[97]^x[67]^x[26]^x[15]^x[3];
	y[2]=x[376]^x[354]^x[339]^x[328]^x[301]^x[290]^x[280]^x[279]^x[274]^x[273]^x[270]^x[269]^x[268]^x[267]^x[263]^x[262]^x[259]^x[258]^x[256]^x[239]^x[238]^x[237]^x[228]^x[226]^x[179]^x[172]^x[168]^x[135]^x[120]^x[119]^x[110]^x[109]^x[108]^x[107]^x[104]^x[99]^x[96]^x[66]^x[25]^x[14]^x[2];
	y[1]=x[375]^x[353]^x[338]^x[327]^x[300]^x[289]^x[279]^x[278]^x[273]^x[272]^x[269]^x[268]^x[267]^x[262]^x[261]^x[258]^x[257]^x[238]^x[237]^x[236]^x[227]^x[225]^x[178]^x[171]^x[167]^x[134]^x[119]^x[118]^x[109]^x[108]^x[107]^x[103]^x[98]^x[65]^x[24]^x[13]^x[1];
	y[0]=x[374]^x[352]^x[337]^x[326]^x[299]^x[288]^x[278]^x[272]^x[268]^x[267]^x[261]^x[257]^x[256]^x[237]^x[236]^x[235]^x[226]^x[224]^x[177]^x[171]^x[166]^x[160]^x[133]^x[118]^x[108]^x[107]^x[102]^x[97]^x[64]^x[23]^x[12]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint53(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[379]^x[378]^x[377]^x[375]^x[374]^x[373]^x[369]^x[367]^x[363]^x[362]^x[358]^x[357]^x[356]^x[353]^x[351]^x[341]^x[331]^x[320]^x[314]^x[313]^x[304]^x[302]^x[293]^x[287]^x[286]^x[277]^x[275]^x[266]^x[253]^x[250]^x[247]^x[246]^x[244]^x[242]^x[240]^x[238]^x[236]^x[235]^x[234]^x[231]^x[229]^x[228]^x[225]^x[223]^x[215]^x[214]^x[213]^x[203]^x[202]^x[193]^x[149]^x[148]^x[147]^x[140]^x[139]^x[129]^x[128]^x[93]^x[90]^x[86]^x[82]^x[78]^x[75]^x[74]^x[72]^x[71]^x[63]^x[57]^x[51]^x[45]^x[17];
	y[30]=x[382]^x[376]^x[374]^x[373]^x[372]^x[368]^x[367]^x[366]^x[362]^x[361]^x[357]^x[356]^x[355]^x[352]^x[351]^x[350]^x[340]^x[286]^x[285]^x[276]^x[274]^x[265]^x[254]^x[252]^x[248]^x[246]^x[245]^x[242]^x[241]^x[239]^x[236]^x[235]^x[234]^x[233]^x[231]^x[230]^x[228]^x[227]^x[225]^x[224]^x[222]^x[214]^x[213]^x[212]^x[202]^x[201]^x[192]^x[158]^x[146]^x[139]^x[138]^x[128]^x[94]^x[92]^x[85]^x[82]^x[81]^x[74]^x[73]^x[71]^x[70]^x[62]^x[56]^x[50]^x[44]^x[16];
	y[29]=x[383]^x[381]^x[377]^x[375]^x[373]^x[372]^x[371]^x[367]^x[366]^x[365]^x[362]^x[361]^x[360]^x[356]^x[355]^x[354]^x[350]^x[349]^x[339]^x[285]^x[284]^x[275]^x[273]^x[264]^x[253]^x[251]^x[247]^x[245]^x[244]^x[241]^x[240]^x[238]^x[234]^x[233]^x[232]^x[230]^x[229]^x[227]^x[226]^x[223]^x[221]^x[213]^x[212]^x[211]^x[202]^x[201]^x[200]^x[159]^x[157]^x[147]^x[145]^x[137]^x[93]^x[91]^x[84]^x[81]^x[80]^x[73]^x[72]^x[70]^x[69]^x[61]^x[55]^x[49]^x[43]^x[15];
	y[28]=x[382]^x[380]^x[376]^x[374]^x[372]^x[371]^x[370]^x[366]^x[365]^x[364]^x[361]^x[360]^x[359]^x[355]^x[354]^x[353]^x[349]^x[348]^x[338]^x[284]^x[283]^x[274]^x[272]^x[263]^x[252]^x[250]^x[246]^x[244]^x[243]^x[240]^x[239]^x[237]^x[233]^x[232]^x[231]^x[229]^x[228]^x[226]^x[225]^x[222]^x[220]^x[212]^x[211]^x[210]^x[201]^x[200]^x[199]^x[158]^x[156]^x[146]^x[144]^x[136]^x[92]^x[90]^x[83]^x[80]^x[79]^x[72]^x[71]^x[69]^x[68]^x[60]^x[54]^x[48]^x[42]^x[14];
	y[27]=x[381]^x[379]^x[375]^x[373]^x[371]^x[370]^x[369]^x[365]^x[364]^x[363]^x[360]^x[359]^x[358]^x[354]^x[353]^x[352]^x[348]^x[347]^x[337]^x[283]^x[282]^x[273]^x[271]^x[262]^x[251]^x[249]^x[245]^x[243]^x[242]^x[239]^x[238]^x[236]^x[232]^x[231]^x[230]^x[228]^x[227]^x[225]^x[224]^x[221]^x[219]^x[211]^x[210]^x[209]^x[200]^x[199]^x[198]^x[157]^x[155]^x[145]^x[143]^x[135]^x[91]^x[89]^x[82]^x[79]^x[78]^x[71]^x[70]^x[68]^x[67]^x[59]^x[53]^x[47]^x[41]^x[13];
	y[26]=x[383]^x[380]^x[378]^x[373]^x[372]^x[370]^x[369]^x[368]^x[364]^x[359]^x[358]^x[357]^x[353]^x[352]^x[347]^x[346]^x[336]^x[319]^x[318]^x[309]^x[308]^x[307]^x[299]^x[288]^x[282]^x[281]^x[272]^x[270]^x[261]^x[253]^x[250]^x[248]^x[245]^x[243]^x[242]^x[241]^x[238]^x[237]^x[235]^x[233]^x[230]^x[229]^x[227]^x[226]^x[224]^x[220]^x[218]^x[210]^x[209]^x[208]^x[199]^x[198]^x[197]^x[156]^x[144]^x[142]^x[134]^x[133]^x[127]^x[106]^x[90]^x[88]^x[85]^x[84]^x[83]^x[81]^x[79]^x[70]^x[69]^x[67]^x[66]^x[58]^x[52]^x[46]^x[40]^x[12];
	y[25]=x[383]^x[382]^x[379]^x[377]^x[373]^x[372]^x[371]^x[369]^x[368]^x[367]^x[363]^x[358]^x[357]^x[356]^x[352]^x[346]^x[345]^x[335]^x[317]^x[308]^x[306]^x[281]^x[280]^x[271]^x[269]^x[260]^x[255]^x[252]^x[249]^x[247]^x[244]^x[242]^x[241]^x[240]^x[237]^x[236]^x[232]^x[229]^x[228]^x[226]^x[225]^x[219]^x[217]^x[209]^x[208]^x[207]^x[198]^x[197]^x[196]^x[155]^x[153]^x[143]^x[141]^x[133]^x[126]^x[105]^x[95]^x[87]^x[84]^x[82]^x[80]^x[78]^x[77]^x[74]^x[69]^x[66]^x[65]^x[57]^x[51]^x[45]^x[39]^x[11];
	y[24]=x[383]^x[382]^x[381]^x[378]^x[376]^x[372]^x[371]^x[370]^x[368]^x[367]^x[366]^x[357]^x[356]^x[355]^x[345]^x[344]^x[334]^x[316]^x[307]^x[305]^x[280]^x[279]^x[270]^x[268]^x[259]^x[254]^x[251]^x[248]^x[246]^x[243]^x[241]^x[240]^x[239]^x[236]^x[235]^x[231]^x[228]^x[227]^x[225]^x[224]^x[218]^x[216]^x[208]^x[207]^x[206]^x[197]^x[196]^x[195]^x[154]^x[152]^x[142]^x[140]^x[132]^x[125]^x[104]^x[94]^x[86]^x[83]^x[81]^x[79]^x[77]^x[76]^x[73]^x[68]^x[65]^x[64]^x[56]^x[50]^x[44]^x[38]^x[10];
	y[23]=x[382]^x[381]^x[380]^x[377]^x[375]^x[371]^x[370]^x[369]^x[367]^x[366]^x[365]^x[356]^x[355]^x[354]^x[344]^x[343]^x[333]^x[315]^x[306]^x[304]^x[279]^x[278]^x[269]^x[267]^x[258]^x[253]^x[250]^x[247]^x[242]^x[240]^x[238]^x[230]^x[228]^x[227]^x[226]^x[217]^x[215]^x[207]^x[206]^x[205]^x[196]^x[195]^x[194]^x[153]^x[151]^x[141]^x[139]^x[131]^x[124]^x[103]^x[93]^x[82]^x[80]^x[78]^x[76]^x[74]^x[72]^x[67]^x[55]^x[49]^x[43]^x[37]^x[9];
	y[22]=x[381]^x[380]^x[379]^x[376]^x[374]^x[370]^x[369]^x[368]^x[366]^x[365]^x[364]^x[355]^x[354]^x[353]^x[343]^x[342]^x[332]^x[314]^x[305]^x[303]^x[278]^x[277]^x[268]^x[266]^x[257]^x[252]^x[249]^x[246]^x[241]^x[239]^x[237]^x[229]^x[227]^x[226]^x[225]^x[216]^x[214]^x[206]^x[205]^x[204]^x[195]^x[194]^x[193]^x[152]^x[150]^x[140]^x[138]^x[130]^x[123]^x[102]^x[92]^x[81]^x[79]^x[77]^x[75]^x[73]^x[71]^x[66]^x[54]^x[48]^x[42]^x[36]^x[8];
	y[21]=x[380]^x[379]^x[378]^x[375]^x[373]^x[369]^x[368]^x[367]^x[365]^x[364]^x[363]^x[354]^x[353]^x[352]^x[342]^x[341]^x[331]^x[313]^x[304]^x[302]^x[277]^x[276]^x[267]^x[265]^x[256]^x[251]^x[248]^x[240]^x[239]^x[238]^x[236]^x[234]^x[226]^x[225]^x[224]^x[215]^x[213]^x[205]^x[204]^x[203]^x[194]^x[193]^x[192]^x[151]^x[149]^x[138]^x[137]^x[129]^x[128]^x[122]^x[101]^x[91]^x[85]^x[80]^x[78]^x[76]^x[72]^x[70]^x[65]^x[53]^x[47]^x[41]^x[35]^x[7];
	y[20]=x[383]^x[379]^x[378]^x[377]^x[374]^x[372]^x[366]^x[364]^x[363]^x[357]^x[353]^x[352]^x[341]^x[340]^x[330]^x[314]^x[313]^x[302]^x[287]^x[276]^x[275]^x[264]^x[255]^x[254]^x[253]^x[250]^x[249]^x[248]^x[247]^x[244]^x[242]^x[238]^x[236]^x[235]^x[234]^x[228]^x[224]^x[223]^x[214]^x[212]^x[204]^x[203]^x[193]^x[192]^x[159]^x[158]^x[150]^x[138]^x[137]^x[136]^x[128]^x[95]^x[94]^x[93]^x[90]^x[82]^x[78]^x[75]^x[74]^x[72]^x[69]^x[64]^x[52]^x[46]^x[40]^x[34]^x[6];
	y[19]=x[383]^x[382]^x[378]^x[377]^x[376]^x[373]^x[371]^x[367]^x[365]^x[363]^x[352]^x[340]^x[339]^x[329]^x[286]^x[275]^x[274]^x[263]^x[255]^x[254]^x[253]^x[252]^x[249]^x[248]^x[247]^x[246]^x[243]^x[241]^x[237]^x[235]^x[233]^x[227]^x[223]^x[222]^x[213]^x[211]^x[203]^x[192]^x[159]^x[157]^x[149]^x[147]^x[138]^x[137]^x[136]^x[135]^x[95]^x[94]^x[93]^x[92]^x[83]^x[81]^x[73]^x[51]^x[45]^x[39]^x[33]^x[5];
	y[18]=x[383]^x[382]^x[381]^x[377]^x[376]^x[375]^x[372]^x[370]^x[366]^x[364]^x[339]^x[338]^x[328]^x[285]^x[274]^x[273]^x[262]^x[254]^x[253]^x[252]^x[251]^x[248]^x[247]^x[246]^x[245]^x[242]^x[240]^x[236]^x[234]^x[232]^x[226]^x[223]^x[222]^x[221]^x[212]^x[210]^x[158]^x[156]^x[148]^x[146]^x[137]^x[136]^x[135]^x[134]^x[94]^x[93]^x[92]^x[91]^x[82]^x[80]^x[72]^x[50]^x[44]^x[38]^x[32]^x[4];
	y[17]=x[382]^x[381]^x[380]^x[376]^x[375]^x[374]^x[371]^x[369]^x[365]^x[363]^x[338]^x[337]^x[327]^x[310]^x[309]^x[298]^x[288]^x[284]^x[273]^x[272]^x[261]^x[253]^x[252]^x[251]^x[250]^x[247]^x[246]^x[245]^x[244]^x[241]^x[239]^x[234]^x[233]^x[231]^x[225]^x[224]^x[222]^x[221]^x[220]^x[211]^x[209]^x[157]^x[155]^x[147]^x[145]^x[136]^x[135]^x[134]^x[133]^x[93]^x[92]^x[91]^x[90]^x[81]^x[79]^x[75]^x[74]^x[71]^x[69]^x[68]^x[64]^x[49]^x[43]^x[37]^x[3];
	y[16]=x[381]^x[380]^x[379]^x[375]^x[374]^x[373]^x[370]^x[368]^x[364]^x[362]^x[337]^x[336]^x[326]^x[308]^x[297]^x[283]^x[272]^x[271]^x[260]^x[252]^x[251]^x[250]^x[249]^x[246]^x[245]^x[244]^x[243]^x[240]^x[238]^x[234]^x[233]^x[232]^x[230]^x[224]^x[221]^x[220]^x[219]^x[210]^x[208]^x[156]^x[154]^x[146]^x[144]^x[135]^x[134]^x[133]^x[132]^x[92]^x[91]^x[90]^x[89]^x[80]^x[78]^x[73]^x[70]^x[67]^x[48]^x[42]^x[36]^x[2];
	y[15]=x[380]^x[379]^x[378]^x[374]^x[373]^x[372]^x[369]^x[367]^x[362]^x[361]^x[352]^x[336]^x[335]^x[325]^x[309]^x[307]^x[298]^x[296]^x[282]^x[271]^x[270]^x[259]^x[251]^x[250]^x[249]^x[248]^x[245]^x[244]^x[243]^x[242]^x[239]^x[237]^x[234]^x[233]^x[232]^x[231]^x[229]^x[220]^x[219]^x[218]^x[209]^x[207]^x[155]^x[153]^x[145]^x[143]^x[134]^x[133]^x[132]^x[131]^x[91]^x[90]^x[89]^x[88]^x[79]^x[77]^x[74]^x[72]^x[69]^x[68]^x[66]^x[47]^x[41]^x[35]^x[1];
	y[14]=x[379]^x[378]^x[377]^x[373]^x[372]^x[371]^x[368]^x[366]^x[362]^x[361]^x[360]^x[335]^x[334]^x[324]^x[308]^x[306]^x[297]^x[295]^x[281]^x[270]^x[269]^x[258]^x[250]^x[249]^x[248]^x[247]^x[244]^x[243]^x[242]^x[241]^x[238]^x[236]^x[233]^x[232]^x[231]^x[230]^x[228]^x[219]^x[218]^x[217]^x[208]^x[206]^x[154]^x[152]^x[144]^x[142]^x[133]^x[132]^x[131]^x[130]^x[90]^x[89]^x[88]^x[87]^x[78]^x[76]^x[73]^x[71]^x[68]^x[67]^x[65]^x[46]^x[40]^x[34]^x[0];
	y[13]=x[378]^x[377]^x[376]^x[372]^x[371]^x[370]^x[367]^x[365]^x[361]^x[360]^x[359]^x[334]^x[333]^x[323]^x[307]^x[305]^x[296]^x[294]^x[280]^x[269]^x[268]^x[257]^x[249]^x[248]^x[247]^x[246]^x[243]^x[242]^x[241]^x[240]^x[237]^x[235]^x[232]^x[231]^x[230]^x[229]^x[227]^x[218]^x[217]^x[216]^x[207]^x[205]^x[153]^x[151]^x[143]^x[141]^x[132]^x[131]^x[130]^x[129]^x[89]^x[88]^x[87]^x[86]^x[77]^x[75]^x[72]^x[70]^x[67]^x[66]^x[64]^x[45]^x[39]^x[33];
	y[12]=x[377]^x[376]^x[375]^x[371]^x[370]^x[369]^x[366]^x[364]^x[360]^x[359]^x[358]^x[333]^x[332]^x[322]^x[306]^x[304]^x[295]^x[293]^x[279]^x[268]^x[267]^x[256]^x[248]^x[247]^x[246]^x[242]^x[241]^x[240]^x[236]^x[231]^x[230]^x[229]^x[226]^x[217]^x[216]^x[215]^x[206]^x[204]^x[152]^x[150]^x[142]^x[140]^x[131]^x[130]^x[129]^x[128]^x[88]^x[87]^x[86]^x[76]^x[71]^x[69]^x[66]^x[65]^x[44]^x[38]^x[32];
	y[11]=x[376]^x[375]^x[374]^x[370]^x[369]^x[368]^x[365]^x[363]^x[359]^x[358]^x[357]^x[332]^x[331]^x[321]^x[305]^x[304]^x[294]^x[293]^x[278]^x[267]^x[247]^x[246]^x[241]^x[240]^x[230]^x[229]^x[225]^x[224]^x[216]^x[215]^x[214]^x[205]^x[203]^x[151]^x[150]^x[141]^x[130]^x[129]^x[128]^x[87]^x[86]^x[70]^x[69]^x[65]^x[43]^x[37];
	y[10]=x[375]^x[374]^x[373]^x[369]^x[368]^x[367]^x[364]^x[362]^x[358]^x[357]^x[356]^x[331]^x[330]^x[320]^x[304]^x[293]^x[277]^x[266]^x[246]^x[245]^x[240]^x[239]^x[234]^x[229]^x[228]^x[224]^x[215]^x[214]^x[213]^x[204]^x[202]^x[150]^x[140]^x[138]^x[129]^x[128]^x[86]^x[85]^x[74]^x[69]^x[64]^x[42]^x[36];
	y[9]=x[378]^x[374]^x[373]^x[372]^x[368]^x[367]^x[366]^x[363]^x[361]^x[357]^x[355]^x[351]^x[329]^x[276]^x[265]^x[255]^x[254]^x[249]^x[248]^x[245]^x[244]^x[243]^x[242]^x[239]^x[238]^x[237]^x[236]^x[234]^x[233]^x[231]^x[228]^x[227]^x[225]^x[214]^x[213]^x[212]^x[203]^x[201]^x[149]^x[148]^x[147]^x[139]^x[137]^x[128]^x[95]^x[94]^x[85]^x[84]^x[83]^x[82]^x[74]^x[73]^x[71]^x[41]^x[35];
	y[8]=x[373]^x[372]^x[371]^x[367]^x[366]^x[365]^x[362]^x[360]^x[356]^x[354]^x[350]^x[328]^x[275]^x[264]^x[254]^x[253]^x[248]^x[247]^x[244]^x[243]^x[242]^x[241]^x[238]^x[237]^x[236]^x[235]^x[233]^x[232]^x[230]^x[227]^x[226]^x[224]^x[213]^x[212]^x[211]^x[202]^x[200]^x[159]^x[148]^x[146]^x[136]^x[94]^x[93]^x[84]^x[83]^x[82]^x[81]^x[73]^x[72]^x[70]^x[40]^x[34];
	y[7]=x[372]^x[371]^x[370]^x[366]^x[365]^x[364]^x[361]^x[359]^x[355]^x[353]^x[349]^x[327]^x[274]^x[263]^x[253]^x[252]^x[247]^x[246]^x[243]^x[242]^x[241]^x[240]^x[237]^x[236]^x[235]^x[232]^x[231]^x[229]^x[226]^x[225]^x[212]^x[211]^x[210]^x[201]^x[199]^x[158]^x[147]^x[145]^x[135]^x[93]^x[92]^x[83]^x[82]^x[81]^x[80]^x[72]^x[71]^x[69]^x[39]^x[33];
	y[6]=x[371]^x[370]^x[369]^x[365]^x[364]^x[363]^x[360]^x[358]^x[354]^x[352]^x[348]^x[326]^x[273]^x[262]^x[252]^x[251]^x[246]^x[245]^x[242]^x[241]^x[240]^x[239]^x[236]^x[235]^x[234]^x[231]^x[230]^x[228]^x[225]^x[224]^x[211]^x[210]^x[209]^x[200]^x[198]^x[157]^x[146]^x[144]^x[134]^x[92]^x[91]^x[82]^x[81]^x[80]^x[79]^x[71]^x[70]^x[68]^x[38]^x[32];
	y[5]=x[374]^x[370]^x[369]^x[368]^x[359]^x[357]^x[352]^x[347]^x[325]^x[310]^x[288]^x[272]^x[261]^x[251]^x[250]^x[245]^x[244]^x[241]^x[240]^x[239]^x[238]^x[234]^x[233]^x[230]^x[229]^x[227]^x[210]^x[209]^x[208]^x[199]^x[197]^x[156]^x[145]^x[143]^x[106]^x[91]^x[90]^x[81]^x[80]^x[79]^x[78]^x[75]^x[70]^x[67]^x[64]^x[37];
	y[4]=x[369]^x[368]^x[367]^x[358]^x[356]^x[346]^x[324]^x[309]^x[298]^x[271]^x[260]^x[250]^x[249]^x[244]^x[243]^x[240]^x[239]^x[238]^x[237]^x[233]^x[232]^x[229]^x[228]^x[226]^x[209]^x[208]^x[207]^x[198]^x[196]^x[155]^x[144]^x[142]^x[132]^x[105]^x[90]^x[89]^x[80]^x[79]^x[78]^x[77]^x[74]^x[69]^x[66]^x[36];
	y[3]=x[368]^x[367]^x[366]^x[357]^x[355]^x[345]^x[323]^x[308]^x[297]^x[270]^x[259]^x[249]^x[248]^x[243]^x[242]^x[239]^x[238]^x[237]^x[236]^x[232]^x[231]^x[228]^x[227]^x[225]^x[208]^x[207]^x[206]^x[197]^x[195]^x[154]^x[143]^x[141]^x[131]^x[104]^x[89]^x[88]^x[79]^x[78]^x[77]^x[76]^x[73]^x[68]^x[65]^x[35];
	y[2]=x[367]^x[366]^x[365]^x[356]^x[354]^x[344]^x[322]^x[307]^x[296]^x[269]^x[258]^x[248]^x[247]^x[242]^x[241]^x[238]^x[237]^x[236]^x[235]^x[231]^x[230]^x[227]^x[226]^x[224]^x[207]^x[206]^x[205]^x[196]^x[194]^x[153]^x[142]^x[140]^x[130]^x[103]^x[88]^x[87]^x[78]^x[77]^x[76]^x[75]^x[72]^x[67]^x[64]^x[34];
	y[1]=x[366]^x[365]^x[364]^x[355]^x[353]^x[343]^x[321]^x[306]^x[295]^x[268]^x[257]^x[247]^x[246]^x[241]^x[240]^x[237]^x[236]^x[235]^x[230]^x[229]^x[226]^x[225]^x[206]^x[205]^x[204]^x[195]^x[193]^x[152]^x[141]^x[139]^x[129]^x[102]^x[87]^x[86]^x[77]^x[76]^x[75]^x[71]^x[66]^x[33];
	y[0]=x[365]^x[364]^x[363]^x[354]^x[352]^x[342]^x[320]^x[305]^x[294]^x[267]^x[256]^x[246]^x[240]^x[236]^x[235]^x[229]^x[225]^x[224]^x[205]^x[204]^x[203]^x[194]^x[192]^x[151]^x[140]^x[139]^x[101]^x[86]^x[76]^x[75]^x[70]^x[65]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint54(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[380]^x[369]^x[351]^x[347]^x[346]^x[345]^x[343]^x[342]^x[341]^x[337]^x[335]^x[331]^x[330]^x[326]^x[325]^x[324]^x[321]^x[319]^x[309]^x[299]^x[288]^x[282]^x[281]^x[272]^x[270]^x[261]^x[255]^x[254]^x[245]^x[243]^x[234]^x[221]^x[218]^x[215]^x[214]^x[212]^x[210]^x[208]^x[206]^x[204]^x[203]^x[202]^x[199]^x[197]^x[196]^x[193]^x[191]^x[183]^x[182]^x[181]^x[171]^x[170]^x[161]^x[145]^x[139]^x[117]^x[116]^x[115]^x[108]^x[107]^x[97]^x[96]^x[61]^x[58]^x[54]^x[50]^x[46]^x[43]^x[42]^x[40]^x[39]^x[31]^x[25]^x[19]^x[13];
	y[30]=x[379]^x[368]^x[350]^x[344]^x[342]^x[341]^x[340]^x[336]^x[335]^x[334]^x[330]^x[329]^x[325]^x[324]^x[323]^x[320]^x[319]^x[318]^x[308]^x[254]^x[253]^x[244]^x[242]^x[233]^x[222]^x[220]^x[216]^x[214]^x[213]^x[210]^x[209]^x[207]^x[204]^x[203]^x[202]^x[201]^x[199]^x[198]^x[196]^x[195]^x[193]^x[192]^x[190]^x[182]^x[181]^x[180]^x[170]^x[169]^x[160]^x[144]^x[138]^x[126]^x[114]^x[107]^x[106]^x[96]^x[62]^x[60]^x[53]^x[50]^x[49]^x[42]^x[41]^x[39]^x[38]^x[30]^x[24]^x[18]^x[12];
	y[29]=x[378]^x[367]^x[351]^x[349]^x[345]^x[343]^x[341]^x[340]^x[339]^x[335]^x[334]^x[333]^x[330]^x[329]^x[328]^x[324]^x[323]^x[322]^x[318]^x[317]^x[307]^x[253]^x[252]^x[243]^x[241]^x[232]^x[221]^x[219]^x[215]^x[213]^x[212]^x[209]^x[208]^x[206]^x[202]^x[201]^x[200]^x[198]^x[197]^x[195]^x[194]^x[191]^x[189]^x[181]^x[180]^x[179]^x[170]^x[169]^x[168]^x[143]^x[137]^x[127]^x[125]^x[115]^x[113]^x[105]^x[61]^x[59]^x[52]^x[49]^x[48]^x[41]^x[40]^x[38]^x[37]^x[29]^x[23]^x[17]^x[11];
	y[28]=x[377]^x[366]^x[350]^x[348]^x[344]^x[342]^x[340]^x[339]^x[338]^x[334]^x[333]^x[332]^x[329]^x[328]^x[327]^x[323]^x[322]^x[321]^x[317]^x[316]^x[306]^x[252]^x[251]^x[242]^x[240]^x[231]^x[220]^x[218]^x[214]^x[212]^x[211]^x[208]^x[207]^x[205]^x[201]^x[200]^x[199]^x[197]^x[196]^x[194]^x[193]^x[190]^x[188]^x[180]^x[179]^x[178]^x[169]^x[168]^x[167]^x[142]^x[136]^x[126]^x[124]^x[114]^x[112]^x[104]^x[60]^x[58]^x[51]^x[48]^x[47]^x[40]^x[39]^x[37]^x[36]^x[28]^x[22]^x[16]^x[10];
	y[27]=x[376]^x[365]^x[349]^x[347]^x[343]^x[341]^x[339]^x[338]^x[337]^x[333]^x[332]^x[331]^x[328]^x[327]^x[326]^x[322]^x[321]^x[320]^x[316]^x[315]^x[305]^x[251]^x[250]^x[241]^x[239]^x[230]^x[219]^x[217]^x[213]^x[211]^x[210]^x[207]^x[206]^x[204]^x[200]^x[199]^x[198]^x[196]^x[195]^x[193]^x[192]^x[189]^x[187]^x[179]^x[178]^x[177]^x[168]^x[167]^x[166]^x[141]^x[135]^x[125]^x[123]^x[113]^x[111]^x[103]^x[59]^x[57]^x[50]^x[47]^x[46]^x[39]^x[38]^x[36]^x[35]^x[27]^x[21]^x[15]^x[9];
	y[26]=x[375]^x[364]^x[351]^x[348]^x[346]^x[341]^x[340]^x[338]^x[337]^x[336]^x[332]^x[327]^x[326]^x[325]^x[321]^x[320]^x[315]^x[314]^x[304]^x[287]^x[286]^x[277]^x[276]^x[275]^x[267]^x[256]^x[250]^x[249]^x[240]^x[238]^x[229]^x[221]^x[218]^x[216]^x[213]^x[211]^x[210]^x[209]^x[206]^x[205]^x[203]^x[201]^x[198]^x[197]^x[195]^x[194]^x[192]^x[188]^x[186]^x[178]^x[177]^x[176]^x[167]^x[166]^x[165]^x[140]^x[134]^x[124]^x[112]^x[110]^x[102]^x[101]^x[95]^x[74]^x[58]^x[56]^x[53]^x[52]^x[51]^x[49]^x[47]^x[38]^x[37]^x[35]^x[34]^x[26]^x[20]^x[14]^x[8];
	y[25]=x[374]^x[363]^x[351]^x[350]^x[347]^x[345]^x[341]^x[340]^x[339]^x[337]^x[336]^x[335]^x[331]^x[326]^x[325]^x[324]^x[320]^x[314]^x[313]^x[303]^x[285]^x[276]^x[274]^x[249]^x[248]^x[239]^x[237]^x[228]^x[223]^x[220]^x[217]^x[215]^x[212]^x[210]^x[209]^x[208]^x[205]^x[204]^x[200]^x[197]^x[196]^x[194]^x[193]^x[187]^x[185]^x[177]^x[176]^x[175]^x[166]^x[165]^x[164]^x[139]^x[133]^x[123]^x[121]^x[111]^x[109]^x[101]^x[94]^x[73]^x[63]^x[55]^x[52]^x[50]^x[48]^x[46]^x[45]^x[42]^x[37]^x[34]^x[33]^x[25]^x[19]^x[13]^x[7];
	y[24]=x[373]^x[362]^x[351]^x[350]^x[349]^x[346]^x[344]^x[340]^x[339]^x[338]^x[336]^x[335]^x[334]^x[325]^x[324]^x[323]^x[313]^x[312]^x[302]^x[284]^x[275]^x[273]^x[248]^x[247]^x[238]^x[236]^x[227]^x[222]^x[219]^x[216]^x[214]^x[211]^x[209]^x[208]^x[207]^x[204]^x[203]^x[199]^x[196]^x[195]^x[193]^x[192]^x[186]^x[184]^x[176]^x[175]^x[174]^x[165]^x[164]^x[163]^x[138]^x[132]^x[122]^x[120]^x[110]^x[108]^x[100]^x[93]^x[72]^x[62]^x[54]^x[51]^x[49]^x[47]^x[45]^x[44]^x[41]^x[36]^x[33]^x[32]^x[24]^x[18]^x[12]^x[6];
	y[23]=x[372]^x[361]^x[350]^x[349]^x[348]^x[345]^x[343]^x[339]^x[338]^x[337]^x[335]^x[334]^x[333]^x[324]^x[323]^x[322]^x[312]^x[311]^x[301]^x[283]^x[274]^x[272]^x[247]^x[246]^x[237]^x[235]^x[226]^x[221]^x[218]^x[215]^x[210]^x[208]^x[206]^x[198]^x[196]^x[195]^x[194]^x[185]^x[183]^x[175]^x[174]^x[173]^x[164]^x[163]^x[162]^x[137]^x[131]^x[121]^x[119]^x[109]^x[107]^x[99]^x[92]^x[71]^x[61]^x[50]^x[48]^x[46]^x[44]^x[42]^x[40]^x[35]^x[23]^x[17]^x[11]^x[5];
	y[22]=x[371]^x[360]^x[349]^x[348]^x[347]^x[344]^x[342]^x[338]^x[337]^x[336]^x[334]^x[333]^x[332]^x[323]^x[322]^x[321]^x[311]^x[310]^x[300]^x[282]^x[273]^x[271]^x[246]^x[245]^x[236]^x[234]^x[225]^x[220]^x[217]^x[214]^x[209]^x[207]^x[205]^x[197]^x[195]^x[194]^x[193]^x[184]^x[182]^x[174]^x[173]^x[172]^x[163]^x[162]^x[161]^x[136]^x[130]^x[120]^x[118]^x[108]^x[106]^x[98]^x[91]^x[70]^x[60]^x[49]^x[47]^x[45]^x[43]^x[41]^x[39]^x[34]^x[22]^x[16]^x[10]^x[4];
	y[21]=x[370]^x[359]^x[348]^x[347]^x[346]^x[343]^x[341]^x[337]^x[336]^x[335]^x[333]^x[332]^x[331]^x[322]^x[321]^x[320]^x[310]^x[309]^x[299]^x[281]^x[272]^x[270]^x[245]^x[244]^x[235]^x[233]^x[224]^x[219]^x[216]^x[208]^x[207]^x[206]^x[204]^x[202]^x[194]^x[193]^x[192]^x[183]^x[181]^x[173]^x[172]^x[171]^x[162]^x[161]^x[160]^x[135]^x[129]^x[119]^x[117]^x[106]^x[105]^x[97]^x[96]^x[90]^x[69]^x[59]^x[53]^x[48]^x[46]^x[44]^x[40]^x[38]^x[33]^x[21]^x[15]^x[9]^x[3];
	y[20]=x[369]^x[358]^x[351]^x[347]^x[346]^x[345]^x[342]^x[340]^x[334]^x[332]^x[331]^x[325]^x[321]^x[320]^x[309]^x[308]^x[298]^x[282]^x[281]^x[270]^x[255]^x[244]^x[243]^x[232]^x[223]^x[222]^x[221]^x[218]^x[217]^x[216]^x[215]^x[212]^x[210]^x[206]^x[204]^x[203]^x[202]^x[196]^x[192]^x[191]^x[182]^x[180]^x[172]^x[171]^x[161]^x[160]^x[134]^x[128]^x[127]^x[126]^x[118]^x[106]^x[105]^x[104]^x[96]^x[63]^x[62]^x[61]^x[58]^x[50]^x[46]^x[43]^x[42]^x[40]^x[37]^x[32]^x[20]^x[14]^x[8]^x[2];
	y[19]=x[368]^x[357]^x[351]^x[350]^x[346]^x[345]^x[344]^x[341]^x[339]^x[335]^x[333]^x[331]^x[320]^x[308]^x[307]^x[297]^x[254]^x[243]^x[242]^x[231]^x[223]^x[222]^x[221]^x[220]^x[217]^x[216]^x[215]^x[214]^x[211]^x[209]^x[205]^x[203]^x[201]^x[195]^x[191]^x[190]^x[181]^x[179]^x[171]^x[160]^x[133]^x[127]^x[125]^x[117]^x[115]^x[106]^x[105]^x[104]^x[103]^x[63]^x[62]^x[61]^x[60]^x[51]^x[49]^x[41]^x[19]^x[13]^x[7]^x[1];
	y[18]=x[367]^x[356]^x[351]^x[350]^x[349]^x[345]^x[344]^x[343]^x[340]^x[338]^x[334]^x[332]^x[307]^x[306]^x[296]^x[253]^x[242]^x[241]^x[230]^x[222]^x[221]^x[220]^x[219]^x[216]^x[215]^x[214]^x[213]^x[210]^x[208]^x[204]^x[202]^x[200]^x[194]^x[191]^x[190]^x[189]^x[180]^x[178]^x[132]^x[126]^x[124]^x[116]^x[114]^x[105]^x[104]^x[103]^x[102]^x[62]^x[61]^x[60]^x[59]^x[50]^x[48]^x[40]^x[18]^x[12]^x[6]^x[0];
	y[17]=x[366]^x[355]^x[350]^x[349]^x[348]^x[344]^x[343]^x[342]^x[339]^x[337]^x[333]^x[331]^x[306]^x[305]^x[295]^x[278]^x[277]^x[266]^x[256]^x[252]^x[241]^x[240]^x[229]^x[221]^x[220]^x[219]^x[218]^x[215]^x[214]^x[213]^x[212]^x[209]^x[207]^x[202]^x[201]^x[199]^x[193]^x[192]^x[190]^x[189]^x[188]^x[179]^x[177]^x[131]^x[125]^x[123]^x[115]^x[113]^x[104]^x[103]^x[102]^x[101]^x[61]^x[60]^x[59]^x[58]^x[49]^x[47]^x[43]^x[42]^x[39]^x[37]^x[36]^x[32]^x[17]^x[11]^x[5];
	y[16]=x[365]^x[354]^x[349]^x[348]^x[347]^x[343]^x[342]^x[341]^x[338]^x[336]^x[332]^x[330]^x[305]^x[304]^x[294]^x[276]^x[265]^x[251]^x[240]^x[239]^x[228]^x[220]^x[219]^x[218]^x[217]^x[214]^x[213]^x[212]^x[211]^x[208]^x[206]^x[202]^x[201]^x[200]^x[198]^x[192]^x[189]^x[188]^x[187]^x[178]^x[176]^x[130]^x[124]^x[122]^x[114]^x[112]^x[103]^x[102]^x[101]^x[100]^x[60]^x[59]^x[58]^x[57]^x[48]^x[46]^x[41]^x[38]^x[35]^x[16]^x[10]^x[4];
	y[15]=x[364]^x[353]^x[348]^x[347]^x[346]^x[342]^x[341]^x[340]^x[337]^x[335]^x[330]^x[329]^x[320]^x[304]^x[303]^x[293]^x[277]^x[275]^x[266]^x[264]^x[250]^x[239]^x[238]^x[227]^x[219]^x[218]^x[217]^x[216]^x[213]^x[212]^x[211]^x[210]^x[207]^x[205]^x[202]^x[201]^x[200]^x[199]^x[197]^x[188]^x[187]^x[186]^x[177]^x[175]^x[129]^x[123]^x[121]^x[113]^x[111]^x[102]^x[101]^x[100]^x[99]^x[59]^x[58]^x[57]^x[56]^x[47]^x[45]^x[42]^x[40]^x[37]^x[36]^x[34]^x[15]^x[9]^x[3];
	y[14]=x[363]^x[352]^x[347]^x[346]^x[345]^x[341]^x[340]^x[339]^x[336]^x[334]^x[330]^x[329]^x[328]^x[303]^x[302]^x[292]^x[276]^x[274]^x[265]^x[263]^x[249]^x[238]^x[237]^x[226]^x[218]^x[217]^x[216]^x[215]^x[212]^x[211]^x[210]^x[209]^x[206]^x[204]^x[201]^x[200]^x[199]^x[198]^x[196]^x[187]^x[186]^x[185]^x[176]^x[174]^x[128]^x[122]^x[120]^x[112]^x[110]^x[101]^x[100]^x[99]^x[98]^x[58]^x[57]^x[56]^x[55]^x[46]^x[44]^x[41]^x[39]^x[36]^x[35]^x[33]^x[14]^x[8]^x[2];
	y[13]=x[346]^x[345]^x[344]^x[340]^x[339]^x[338]^x[335]^x[333]^x[329]^x[328]^x[327]^x[302]^x[301]^x[291]^x[275]^x[273]^x[264]^x[262]^x[248]^x[237]^x[236]^x[225]^x[217]^x[216]^x[215]^x[214]^x[211]^x[210]^x[209]^x[208]^x[205]^x[203]^x[200]^x[199]^x[198]^x[197]^x[195]^x[186]^x[185]^x[184]^x[175]^x[173]^x[121]^x[119]^x[111]^x[109]^x[100]^x[99]^x[98]^x[97]^x[57]^x[56]^x[55]^x[54]^x[45]^x[43]^x[40]^x[38]^x[35]^x[34]^x[32]^x[13]^x[7]^x[1];
	y[12]=x[345]^x[344]^x[343]^x[339]^x[338]^x[337]^x[334]^x[332]^x[328]^x[327]^x[326]^x[301]^x[300]^x[290]^x[274]^x[272]^x[263]^x[261]^x[247]^x[236]^x[235]^x[224]^x[216]^x[215]^x[214]^x[210]^x[209]^x[208]^x[204]^x[199]^x[198]^x[197]^x[194]^x[185]^x[184]^x[183]^x[174]^x[172]^x[120]^x[118]^x[110]^x[108]^x[99]^x[98]^x[97]^x[96]^x[56]^x[55]^x[54]^x[44]^x[39]^x[37]^x[34]^x[33]^x[12]^x[6]^x[0];
	y[11]=x[344]^x[343]^x[342]^x[338]^x[337]^x[336]^x[333]^x[331]^x[327]^x[326]^x[325]^x[300]^x[299]^x[289]^x[273]^x[272]^x[262]^x[261]^x[246]^x[235]^x[215]^x[214]^x[209]^x[208]^x[198]^x[197]^x[193]^x[192]^x[184]^x[183]^x[182]^x[173]^x[171]^x[119]^x[118]^x[109]^x[98]^x[97]^x[96]^x[55]^x[54]^x[38]^x[37]^x[33]^x[11]^x[5];
	y[10]=x[343]^x[342]^x[341]^x[337]^x[336]^x[335]^x[332]^x[330]^x[326]^x[325]^x[324]^x[299]^x[298]^x[288]^x[272]^x[261]^x[245]^x[234]^x[214]^x[213]^x[208]^x[207]^x[202]^x[197]^x[196]^x[192]^x[183]^x[182]^x[181]^x[172]^x[170]^x[118]^x[108]^x[106]^x[97]^x[96]^x[54]^x[53]^x[42]^x[37]^x[32]^x[10]^x[4];
	y[9]=x[346]^x[342]^x[341]^x[340]^x[336]^x[335]^x[334]^x[331]^x[329]^x[325]^x[323]^x[319]^x[297]^x[244]^x[233]^x[223]^x[222]^x[217]^x[216]^x[213]^x[212]^x[211]^x[210]^x[207]^x[206]^x[205]^x[204]^x[202]^x[201]^x[199]^x[196]^x[195]^x[193]^x[182]^x[181]^x[180]^x[171]^x[169]^x[117]^x[116]^x[115]^x[107]^x[105]^x[96]^x[63]^x[62]^x[53]^x[52]^x[51]^x[50]^x[42]^x[41]^x[39]^x[9]^x[3];
	y[8]=x[341]^x[340]^x[339]^x[335]^x[334]^x[333]^x[330]^x[328]^x[324]^x[322]^x[318]^x[296]^x[243]^x[232]^x[222]^x[221]^x[216]^x[215]^x[212]^x[211]^x[210]^x[209]^x[206]^x[205]^x[204]^x[203]^x[201]^x[200]^x[198]^x[195]^x[194]^x[192]^x[181]^x[180]^x[179]^x[170]^x[168]^x[127]^x[116]^x[114]^x[104]^x[62]^x[61]^x[52]^x[51]^x[50]^x[49]^x[41]^x[40]^x[38]^x[8]^x[2];
	y[7]=x[340]^x[339]^x[338]^x[334]^x[333]^x[332]^x[329]^x[327]^x[323]^x[321]^x[317]^x[295]^x[242]^x[231]^x[221]^x[220]^x[215]^x[214]^x[211]^x[210]^x[209]^x[208]^x[205]^x[204]^x[203]^x[200]^x[199]^x[197]^x[194]^x[193]^x[180]^x[179]^x[178]^x[169]^x[167]^x[126]^x[115]^x[113]^x[103]^x[61]^x[60]^x[51]^x[50]^x[49]^x[48]^x[40]^x[39]^x[37]^x[7]^x[1];
	y[6]=x[339]^x[338]^x[337]^x[333]^x[332]^x[331]^x[328]^x[326]^x[322]^x[320]^x[316]^x[294]^x[241]^x[230]^x[220]^x[219]^x[214]^x[213]^x[210]^x[209]^x[208]^x[207]^x[204]^x[203]^x[202]^x[199]^x[198]^x[196]^x[193]^x[192]^x[179]^x[178]^x[177]^x[168]^x[166]^x[125]^x[114]^x[112]^x[102]^x[60]^x[59]^x[50]^x[49]^x[48]^x[47]^x[39]^x[38]^x[36]^x[6]^x[0];
	y[5]=x[342]^x[338]^x[337]^x[336]^x[327]^x[325]^x[320]^x[315]^x[293]^x[278]^x[256]^x[240]^x[229]^x[219]^x[218]^x[213]^x[212]^x[209]^x[208]^x[207]^x[206]^x[202]^x[201]^x[198]^x[197]^x[195]^x[178]^x[177]^x[176]^x[167]^x[165]^x[124]^x[113]^x[111]^x[74]^x[59]^x[58]^x[49]^x[48]^x[47]^x[46]^x[43]^x[38]^x[35]^x[32]^x[5];
	y[4]=x[337]^x[336]^x[335]^x[326]^x[324]^x[314]^x[292]^x[277]^x[266]^x[239]^x[228]^x[218]^x[217]^x[212]^x[211]^x[208]^x[207]^x[206]^x[205]^x[201]^x[200]^x[197]^x[196]^x[194]^x[177]^x[176]^x[175]^x[166]^x[164]^x[123]^x[112]^x[110]^x[100]^x[73]^x[58]^x[57]^x[48]^x[47]^x[46]^x[45]^x[42]^x[37]^x[34]^x[4];
	y[3]=x[336]^x[335]^x[334]^x[325]^x[323]^x[313]^x[291]^x[276]^x[265]^x[238]^x[227]^x[217]^x[216]^x[211]^x[210]^x[207]^x[206]^x[205]^x[204]^x[200]^x[199]^x[196]^x[195]^x[193]^x[176]^x[175]^x[174]^x[165]^x[163]^x[122]^x[111]^x[109]^x[99]^x[72]^x[57]^x[56]^x[47]^x[46]^x[45]^x[44]^x[41]^x[36]^x[33]^x[3];
	y[2]=x[335]^x[334]^x[333]^x[324]^x[322]^x[312]^x[290]^x[275]^x[264]^x[237]^x[226]^x[216]^x[215]^x[210]^x[209]^x[206]^x[205]^x[204]^x[203]^x[199]^x[198]^x[195]^x[194]^x[192]^x[175]^x[174]^x[173]^x[164]^x[162]^x[121]^x[110]^x[108]^x[98]^x[71]^x[56]^x[55]^x[46]^x[45]^x[44]^x[43]^x[40]^x[35]^x[32]^x[2];
	y[1]=x[334]^x[333]^x[332]^x[323]^x[321]^x[311]^x[289]^x[274]^x[263]^x[236]^x[225]^x[215]^x[214]^x[209]^x[208]^x[205]^x[204]^x[203]^x[198]^x[197]^x[194]^x[193]^x[174]^x[173]^x[172]^x[163]^x[161]^x[120]^x[109]^x[107]^x[97]^x[70]^x[55]^x[54]^x[45]^x[44]^x[43]^x[39]^x[34]^x[1];
	y[0]=x[333]^x[332]^x[331]^x[322]^x[320]^x[310]^x[288]^x[273]^x[262]^x[235]^x[224]^x[214]^x[208]^x[204]^x[203]^x[197]^x[193]^x[192]^x[173]^x[172]^x[171]^x[162]^x[160]^x[119]^x[108]^x[107]^x[69]^x[54]^x[44]^x[43]^x[38]^x[33]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint55(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[377]^x[376]^x[373]^x[371]^x[367]^x[365]^x[362]^x[356]^x[348]^x[337]^x[319]^x[315]^x[314]^x[313]^x[311]^x[310]^x[309]^x[305]^x[303]^x[299]^x[298]^x[294]^x[293]^x[292]^x[289]^x[287]^x[277]^x[267]^x[256]^x[250]^x[249]^x[240]^x[238]^x[229]^x[223]^x[222]^x[213]^x[211]^x[202]^x[189]^x[186]^x[183]^x[182]^x[180]^x[178]^x[176]^x[174]^x[172]^x[171]^x[170]^x[167]^x[165]^x[164]^x[161]^x[151]^x[150]^x[149]^x[139]^x[138]^x[135]^x[129]^x[113]^x[107]^x[85]^x[84]^x[83]^x[76]^x[75]^x[65]^x[64]^x[29]^x[26]^x[22]^x[18]^x[14]^x[11]^x[10]^x[8]^x[7];
	y[30]=x[382]^x[381]^x[376]^x[375]^x[372]^x[370]^x[366]^x[364]^x[361]^x[355]^x[347]^x[336]^x[318]^x[312]^x[310]^x[309]^x[308]^x[304]^x[303]^x[302]^x[298]^x[297]^x[293]^x[292]^x[291]^x[288]^x[287]^x[286]^x[276]^x[222]^x[221]^x[212]^x[210]^x[201]^x[190]^x[188]^x[184]^x[182]^x[181]^x[178]^x[177]^x[175]^x[172]^x[171]^x[170]^x[169]^x[167]^x[166]^x[164]^x[163]^x[161]^x[160]^x[150]^x[149]^x[148]^x[138]^x[137]^x[134]^x[128]^x[112]^x[106]^x[94]^x[82]^x[75]^x[74]^x[64]^x[30]^x[28]^x[21]^x[18]^x[17]^x[10]^x[9]^x[7]^x[6];
	y[29]=x[381]^x[380]^x[375]^x[374]^x[371]^x[369]^x[365]^x[363]^x[360]^x[354]^x[346]^x[335]^x[319]^x[317]^x[313]^x[311]^x[309]^x[308]^x[307]^x[303]^x[302]^x[301]^x[298]^x[297]^x[296]^x[292]^x[291]^x[290]^x[286]^x[285]^x[275]^x[221]^x[220]^x[211]^x[209]^x[200]^x[189]^x[187]^x[183]^x[181]^x[180]^x[177]^x[176]^x[174]^x[170]^x[169]^x[168]^x[166]^x[165]^x[163]^x[162]^x[159]^x[149]^x[148]^x[147]^x[138]^x[137]^x[136]^x[133]^x[111]^x[105]^x[95]^x[93]^x[83]^x[81]^x[73]^x[29]^x[27]^x[20]^x[17]^x[16]^x[9]^x[8]^x[6]^x[5];
	y[28]=x[380]^x[379]^x[374]^x[373]^x[370]^x[368]^x[364]^x[362]^x[359]^x[353]^x[345]^x[334]^x[318]^x[316]^x[312]^x[310]^x[308]^x[307]^x[306]^x[302]^x[301]^x[300]^x[297]^x[296]^x[295]^x[291]^x[290]^x[289]^x[285]^x[284]^x[274]^x[220]^x[219]^x[210]^x[208]^x[199]^x[188]^x[186]^x[182]^x[180]^x[179]^x[176]^x[175]^x[173]^x[169]^x[168]^x[167]^x[165]^x[164]^x[162]^x[161]^x[158]^x[148]^x[147]^x[146]^x[137]^x[136]^x[135]^x[132]^x[110]^x[104]^x[94]^x[92]^x[82]^x[80]^x[72]^x[28]^x[26]^x[19]^x[16]^x[15]^x[8]^x[7]^x[5]^x[4];
	y[27]=x[379]^x[378]^x[373]^x[372]^x[369]^x[367]^x[363]^x[361]^x[358]^x[352]^x[344]^x[333]^x[317]^x[315]^x[311]^x[309]^x[307]^x[306]^x[305]^x[301]^x[300]^x[299]^x[296]^x[295]^x[294]^x[290]^x[289]^x[288]^x[284]^x[283]^x[273]^x[219]^x[218]^x[209]^x[207]^x[198]^x[187]^x[185]^x[181]^x[179]^x[178]^x[175]^x[174]^x[172]^x[168]^x[167]^x[166]^x[164]^x[163]^x[161]^x[160]^x[157]^x[147]^x[146]^x[145]^x[136]^x[135]^x[134]^x[131]^x[109]^x[103]^x[93]^x[91]^x[81]^x[79]^x[71]^x[27]^x[25]^x[18]^x[15]^x[14]^x[7]^x[6]^x[4]^x[3];
	y[26]=x[383]^x[378]^x[377]^x[372]^x[371]^x[368]^x[366]^x[360]^x[357]^x[343]^x[332]^x[319]^x[316]^x[314]^x[309]^x[308]^x[306]^x[305]^x[304]^x[300]^x[295]^x[294]^x[293]^x[289]^x[288]^x[283]^x[282]^x[272]^x[255]^x[254]^x[245]^x[244]^x[243]^x[235]^x[224]^x[218]^x[217]^x[208]^x[206]^x[197]^x[189]^x[186]^x[184]^x[181]^x[179]^x[178]^x[177]^x[174]^x[173]^x[171]^x[169]^x[166]^x[165]^x[163]^x[162]^x[160]^x[156]^x[146]^x[145]^x[144]^x[135]^x[134]^x[133]^x[130]^x[108]^x[102]^x[92]^x[80]^x[78]^x[70]^x[69]^x[63]^x[42]^x[26]^x[24]^x[21]^x[20]^x[19]^x[17]^x[15]^x[6]^x[5]^x[3]^x[2];
	y[25]=x[382]^x[377]^x[376]^x[371]^x[370]^x[367]^x[365]^x[359]^x[356]^x[342]^x[331]^x[319]^x[318]^x[315]^x[313]^x[309]^x[308]^x[307]^x[305]^x[304]^x[303]^x[299]^x[294]^x[293]^x[292]^x[288]^x[282]^x[281]^x[271]^x[253]^x[244]^x[242]^x[217]^x[216]^x[207]^x[205]^x[196]^x[191]^x[188]^x[185]^x[183]^x[180]^x[178]^x[177]^x[176]^x[173]^x[172]^x[168]^x[165]^x[164]^x[162]^x[161]^x[155]^x[145]^x[144]^x[143]^x[134]^x[133]^x[132]^x[129]^x[107]^x[101]^x[91]^x[89]^x[79]^x[77]^x[69]^x[62]^x[41]^x[31]^x[23]^x[20]^x[18]^x[16]^x[14]^x[13]^x[10]^x[5]^x[2]^x[1];
	y[24]=x[381]^x[376]^x[375]^x[370]^x[369]^x[366]^x[364]^x[358]^x[355]^x[341]^x[330]^x[319]^x[318]^x[317]^x[314]^x[312]^x[308]^x[307]^x[306]^x[304]^x[303]^x[302]^x[293]^x[292]^x[291]^x[281]^x[280]^x[270]^x[252]^x[243]^x[241]^x[216]^x[215]^x[206]^x[204]^x[195]^x[190]^x[187]^x[184]^x[182]^x[179]^x[177]^x[176]^x[175]^x[172]^x[171]^x[167]^x[164]^x[163]^x[161]^x[160]^x[154]^x[144]^x[143]^x[142]^x[133]^x[132]^x[131]^x[128]^x[106]^x[100]^x[90]^x[88]^x[78]^x[76]^x[68]^x[61]^x[40]^x[30]^x[22]^x[19]^x[17]^x[15]^x[13]^x[12]^x[9]^x[4]^x[1]^x[0];
	y[23]=x[380]^x[375]^x[374]^x[369]^x[368]^x[365]^x[363]^x[357]^x[354]^x[340]^x[329]^x[318]^x[317]^x[316]^x[313]^x[311]^x[307]^x[306]^x[305]^x[303]^x[302]^x[301]^x[292]^x[291]^x[290]^x[280]^x[279]^x[269]^x[251]^x[242]^x[240]^x[215]^x[214]^x[205]^x[203]^x[194]^x[189]^x[186]^x[183]^x[178]^x[176]^x[174]^x[166]^x[164]^x[163]^x[162]^x[153]^x[143]^x[142]^x[141]^x[132]^x[131]^x[130]^x[105]^x[99]^x[89]^x[87]^x[77]^x[75]^x[67]^x[60]^x[39]^x[29]^x[18]^x[16]^x[14]^x[12]^x[10]^x[8]^x[3];
	y[22]=x[379]^x[374]^x[373]^x[368]^x[367]^x[364]^x[362]^x[356]^x[353]^x[339]^x[328]^x[317]^x[316]^x[315]^x[312]^x[310]^x[306]^x[305]^x[304]^x[302]^x[301]^x[300]^x[291]^x[290]^x[289]^x[279]^x[278]^x[268]^x[250]^x[241]^x[239]^x[214]^x[213]^x[204]^x[202]^x[193]^x[188]^x[185]^x[182]^x[177]^x[175]^x[173]^x[165]^x[163]^x[162]^x[161]^x[152]^x[142]^x[141]^x[140]^x[131]^x[130]^x[129]^x[104]^x[98]^x[88]^x[86]^x[76]^x[74]^x[66]^x[59]^x[38]^x[28]^x[17]^x[15]^x[13]^x[11]^x[9]^x[7]^x[2];
	y[21]=x[378]^x[373]^x[372]^x[367]^x[366]^x[363]^x[361]^x[355]^x[352]^x[338]^x[327]^x[316]^x[315]^x[314]^x[311]^x[309]^x[305]^x[304]^x[303]^x[301]^x[300]^x[299]^x[290]^x[289]^x[288]^x[278]^x[277]^x[267]^x[249]^x[240]^x[238]^x[213]^x[212]^x[203]^x[201]^x[192]^x[187]^x[184]^x[176]^x[175]^x[174]^x[172]^x[170]^x[162]^x[161]^x[160]^x[151]^x[141]^x[140]^x[139]^x[130]^x[129]^x[128]^x[103]^x[97]^x[87]^x[85]^x[74]^x[73]^x[65]^x[64]^x[58]^x[37]^x[27]^x[21]^x[16]^x[14]^x[12]^x[8]^x[6]^x[1];
	y[20]=x[383]^x[377]^x[372]^x[371]^x[366]^x[365]^x[360]^x[354]^x[337]^x[326]^x[319]^x[315]^x[314]^x[313]^x[310]^x[308]^x[302]^x[300]^x[299]^x[293]^x[289]^x[288]^x[277]^x[276]^x[266]^x[250]^x[249]^x[238]^x[223]^x[212]^x[211]^x[200]^x[191]^x[190]^x[189]^x[186]^x[185]^x[184]^x[183]^x[180]^x[178]^x[174]^x[172]^x[171]^x[170]^x[164]^x[160]^x[159]^x[150]^x[140]^x[139]^x[129]^x[128]^x[102]^x[96]^x[95]^x[94]^x[86]^x[74]^x[73]^x[72]^x[64]^x[31]^x[30]^x[29]^x[26]^x[18]^x[14]^x[11]^x[10]^x[8]^x[5]^x[0];
	y[19]=x[382]^x[376]^x[371]^x[370]^x[365]^x[364]^x[359]^x[353]^x[336]^x[325]^x[319]^x[318]^x[314]^x[313]^x[312]^x[309]^x[307]^x[303]^x[301]^x[299]^x[288]^x[276]^x[275]^x[265]^x[222]^x[211]^x[210]^x[199]^x[191]^x[190]^x[189]^x[188]^x[185]^x[184]^x[183]^x[182]^x[179]^x[177]^x[173]^x[171]^x[169]^x[163]^x[159]^x[158]^x[149]^x[139]^x[128]^x[101]^x[95]^x[93]^x[85]^x[83]^x[74]^x[73]^x[72]^x[71]^x[31]^x[30]^x[29]^x[28]^x[19]^x[17]^x[9];
	y[18]=x[381]^x[375]^x[370]^x[369]^x[364]^x[363]^x[358]^x[352]^x[335]^x[324]^x[319]^x[318]^x[317]^x[313]^x[312]^x[311]^x[308]^x[306]^x[302]^x[300]^x[275]^x[274]^x[264]^x[221]^x[210]^x[209]^x[198]^x[190]^x[189]^x[188]^x[187]^x[184]^x[183]^x[182]^x[181]^x[178]^x[176]^x[172]^x[170]^x[168]^x[162]^x[159]^x[158]^x[157]^x[148]^x[100]^x[94]^x[92]^x[84]^x[82]^x[73]^x[72]^x[71]^x[70]^x[30]^x[29]^x[28]^x[27]^x[18]^x[16]^x[8];
	y[17]=x[380]^x[374]^x[369]^x[368]^x[363]^x[357]^x[334]^x[323]^x[318]^x[317]^x[316]^x[312]^x[311]^x[310]^x[307]^x[305]^x[301]^x[299]^x[274]^x[273]^x[263]^x[246]^x[245]^x[234]^x[224]^x[220]^x[209]^x[208]^x[197]^x[189]^x[188]^x[187]^x[186]^x[183]^x[182]^x[181]^x[180]^x[177]^x[175]^x[170]^x[169]^x[167]^x[161]^x[160]^x[158]^x[157]^x[156]^x[147]^x[99]^x[93]^x[91]^x[83]^x[81]^x[72]^x[71]^x[70]^x[69]^x[29]^x[28]^x[27]^x[26]^x[17]^x[15]^x[11]^x[10]^x[7]^x[5]^x[4]^x[0];
	y[16]=x[379]^x[373]^x[368]^x[367]^x[362]^x[356]^x[333]^x[322]^x[317]^x[316]^x[315]^x[311]^x[310]^x[309]^x[306]^x[304]^x[300]^x[298]^x[273]^x[272]^x[262]^x[244]^x[233]^x[219]^x[208]^x[207]^x[196]^x[188]^x[187]^x[186]^x[185]^x[182]^x[181]^x[180]^x[179]^x[176]^x[174]^x[170]^x[169]^x[168]^x[166]^x[160]^x[157]^x[156]^x[155]^x[146]^x[98]^x[92]^x[90]^x[82]^x[80]^x[71]^x[70]^x[69]^x[68]^x[28]^x[27]^x[26]^x[25]^x[16]^x[14]^x[9]^x[6]^x[3];
	y[15]=x[378]^x[372]^x[367]^x[366]^x[361]^x[355]^x[332]^x[321]^x[316]^x[315]^x[314]^x[310]^x[309]^x[308]^x[305]^x[303]^x[298]^x[297]^x[288]^x[272]^x[271]^x[261]^x[245]^x[243]^x[234]^x[232]^x[218]^x[207]^x[206]^x[195]^x[187]^x[186]^x[185]^x[184]^x[181]^x[180]^x[179]^x[178]^x[175]^x[173]^x[170]^x[169]^x[168]^x[167]^x[165]^x[156]^x[155]^x[154]^x[145]^x[97]^x[91]^x[89]^x[81]^x[79]^x[70]^x[69]^x[68]^x[67]^x[27]^x[26]^x[25]^x[24]^x[15]^x[13]^x[10]^x[8]^x[5]^x[4]^x[2];
	y[14]=x[377]^x[371]^x[366]^x[365]^x[360]^x[354]^x[331]^x[320]^x[315]^x[314]^x[313]^x[309]^x[308]^x[307]^x[304]^x[302]^x[298]^x[297]^x[296]^x[271]^x[270]^x[260]^x[244]^x[242]^x[233]^x[231]^x[217]^x[206]^x[205]^x[194]^x[186]^x[185]^x[184]^x[183]^x[180]^x[179]^x[178]^x[177]^x[174]^x[172]^x[169]^x[168]^x[167]^x[166]^x[164]^x[155]^x[154]^x[153]^x[144]^x[96]^x[90]^x[88]^x[80]^x[78]^x[69]^x[68]^x[67]^x[66]^x[26]^x[25]^x[24]^x[23]^x[14]^x[12]^x[9]^x[7]^x[4]^x[3]^x[1];
	y[13]=x[376]^x[370]^x[365]^x[364]^x[359]^x[353]^x[314]^x[313]^x[312]^x[308]^x[307]^x[306]^x[303]^x[301]^x[297]^x[296]^x[295]^x[270]^x[269]^x[259]^x[243]^x[241]^x[232]^x[230]^x[216]^x[205]^x[204]^x[193]^x[185]^x[184]^x[183]^x[182]^x[179]^x[178]^x[177]^x[176]^x[173]^x[171]^x[168]^x[167]^x[166]^x[165]^x[163]^x[154]^x[153]^x[152]^x[143]^x[89]^x[87]^x[79]^x[77]^x[68]^x[67]^x[66]^x[65]^x[25]^x[24]^x[23]^x[22]^x[13]^x[11]^x[8]^x[6]^x[3]^x[2]^x[0];
	y[12]=x[375]^x[369]^x[364]^x[363]^x[358]^x[352]^x[313]^x[312]^x[311]^x[307]^x[306]^x[305]^x[302]^x[300]^x[296]^x[295]^x[294]^x[269]^x[268]^x[258]^x[242]^x[240]^x[231]^x[229]^x[215]^x[204]^x[203]^x[192]^x[184]^x[183]^x[182]^x[178]^x[177]^x[176]^x[172]^x[167]^x[166]^x[165]^x[162]^x[153]^x[152]^x[151]^x[142]^x[88]^x[86]^x[78]^x[76]^x[67]^x[66]^x[65]^x[64]^x[24]^x[23]^x[22]^x[12]^x[7]^x[5]^x[2]^x[1];
	y[11]=x[374]^x[368]^x[363]^x[357]^x[312]^x[311]^x[310]^x[306]^x[305]^x[304]^x[301]^x[299]^x[295]^x[294]^x[293]^x[268]^x[267]^x[257]^x[241]^x[240]^x[230]^x[229]^x[214]^x[203]^x[183]^x[182]^x[177]^x[176]^x[166]^x[165]^x[161]^x[160]^x[152]^x[151]^x[150]^x[141]^x[87]^x[86]^x[77]^x[66]^x[65]^x[64]^x[23]^x[22]^x[6]^x[5]^x[1];
	y[10]=x[373]^x[367]^x[362]^x[356]^x[311]^x[310]^x[309]^x[305]^x[304]^x[303]^x[300]^x[298]^x[294]^x[293]^x[292]^x[267]^x[266]^x[256]^x[240]^x[229]^x[213]^x[202]^x[182]^x[181]^x[176]^x[175]^x[170]^x[165]^x[164]^x[160]^x[151]^x[150]^x[149]^x[140]^x[86]^x[76]^x[74]^x[65]^x[64]^x[22]^x[21]^x[10]^x[5]^x[0];
	y[9]=x[372]^x[366]^x[361]^x[355]^x[314]^x[310]^x[309]^x[308]^x[304]^x[303]^x[302]^x[299]^x[297]^x[293]^x[291]^x[287]^x[265]^x[212]^x[201]^x[191]^x[190]^x[185]^x[184]^x[181]^x[180]^x[179]^x[178]^x[175]^x[174]^x[173]^x[172]^x[170]^x[169]^x[167]^x[164]^x[163]^x[161]^x[150]^x[149]^x[148]^x[139]^x[85]^x[84]^x[83]^x[75]^x[73]^x[64]^x[31]^x[30]^x[21]^x[20]^x[19]^x[18]^x[10]^x[9]^x[7];
	y[8]=x[371]^x[365]^x[360]^x[354]^x[309]^x[308]^x[307]^x[303]^x[302]^x[301]^x[298]^x[296]^x[292]^x[290]^x[286]^x[264]^x[211]^x[200]^x[190]^x[189]^x[184]^x[183]^x[180]^x[179]^x[178]^x[177]^x[174]^x[173]^x[172]^x[171]^x[169]^x[168]^x[166]^x[163]^x[162]^x[160]^x[149]^x[148]^x[147]^x[138]^x[95]^x[84]^x[82]^x[72]^x[30]^x[29]^x[20]^x[19]^x[18]^x[17]^x[9]^x[8]^x[6];
	y[7]=x[370]^x[364]^x[359]^x[353]^x[308]^x[307]^x[306]^x[302]^x[301]^x[300]^x[297]^x[295]^x[291]^x[289]^x[285]^x[263]^x[210]^x[199]^x[189]^x[188]^x[183]^x[182]^x[179]^x[178]^x[177]^x[176]^x[173]^x[172]^x[171]^x[168]^x[167]^x[165]^x[162]^x[161]^x[148]^x[147]^x[146]^x[137]^x[94]^x[83]^x[81]^x[71]^x[29]^x[28]^x[19]^x[18]^x[17]^x[16]^x[8]^x[7]^x[5];
	y[6]=x[369]^x[363]^x[358]^x[352]^x[307]^x[306]^x[305]^x[301]^x[300]^x[299]^x[296]^x[294]^x[290]^x[288]^x[284]^x[262]^x[209]^x[198]^x[188]^x[187]^x[182]^x[181]^x[178]^x[177]^x[176]^x[175]^x[172]^x[171]^x[170]^x[167]^x[166]^x[164]^x[161]^x[160]^x[147]^x[146]^x[145]^x[136]^x[93]^x[82]^x[80]^x[70]^x[28]^x[27]^x[18]^x[17]^x[16]^x[15]^x[7]^x[6]^x[4];
	y[5]=x[368]^x[357]^x[310]^x[306]^x[305]^x[304]^x[295]^x[293]^x[288]^x[283]^x[261]^x[246]^x[224]^x[208]^x[197]^x[187]^x[186]^x[181]^x[180]^x[177]^x[176]^x[175]^x[174]^x[170]^x[169]^x[166]^x[165]^x[163]^x[146]^x[145]^x[144]^x[135]^x[92]^x[81]^x[79]^x[42]^x[27]^x[26]^x[17]^x[16]^x[15]^x[14]^x[11]^x[6]^x[3]^x[0];
	y[4]=x[367]^x[356]^x[305]^x[304]^x[303]^x[294]^x[292]^x[282]^x[260]^x[245]^x[234]^x[207]^x[196]^x[186]^x[185]^x[180]^x[179]^x[176]^x[175]^x[174]^x[173]^x[169]^x[168]^x[165]^x[164]^x[162]^x[145]^x[144]^x[143]^x[134]^x[91]^x[80]^x[78]^x[68]^x[41]^x[26]^x[25]^x[16]^x[15]^x[14]^x[13]^x[10]^x[5]^x[2];
	y[3]=x[366]^x[355]^x[304]^x[303]^x[302]^x[293]^x[291]^x[281]^x[259]^x[244]^x[233]^x[206]^x[195]^x[185]^x[184]^x[179]^x[178]^x[175]^x[174]^x[173]^x[172]^x[168]^x[167]^x[164]^x[163]^x[161]^x[144]^x[143]^x[142]^x[133]^x[90]^x[79]^x[77]^x[67]^x[40]^x[25]^x[24]^x[15]^x[14]^x[13]^x[12]^x[9]^x[4]^x[1];
	y[2]=x[365]^x[354]^x[303]^x[302]^x[301]^x[292]^x[290]^x[280]^x[258]^x[243]^x[232]^x[205]^x[194]^x[184]^x[183]^x[178]^x[177]^x[174]^x[173]^x[172]^x[171]^x[167]^x[166]^x[163]^x[162]^x[160]^x[143]^x[142]^x[141]^x[132]^x[89]^x[78]^x[76]^x[66]^x[39]^x[24]^x[23]^x[14]^x[13]^x[12]^x[11]^x[8]^x[3]^x[0];
	y[1]=x[364]^x[353]^x[302]^x[301]^x[300]^x[291]^x[289]^x[279]^x[257]^x[242]^x[231]^x[204]^x[193]^x[183]^x[182]^x[177]^x[176]^x[173]^x[172]^x[171]^x[166]^x[165]^x[162]^x[161]^x[142]^x[141]^x[140]^x[131]^x[88]^x[77]^x[75]^x[65]^x[38]^x[23]^x[22]^x[13]^x[12]^x[11]^x[7]^x[2];
	y[0]=x[363]^x[352]^x[301]^x[300]^x[299]^x[290]^x[288]^x[278]^x[256]^x[241]^x[230]^x[203]^x[192]^x[182]^x[176]^x[172]^x[171]^x[165]^x[161]^x[160]^x[141]^x[140]^x[139]^x[130]^x[87]^x[76]^x[75]^x[37]^x[22]^x[12]^x[11]^x[6]^x[1];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint56(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[378]^x[377]^x[373]^x[368]^x[366]^x[364]^x[363]^x[362]^x[359]^x[357]^x[353]^x[351]^x[350]^x[345]^x[344]^x[341]^x[339]^x[335]^x[333]^x[330]^x[324]^x[316]^x[305]^x[287]^x[283]^x[282]^x[281]^x[279]^x[278]^x[277]^x[273]^x[271]^x[267]^x[266]^x[262]^x[261]^x[260]^x[257]^x[255]^x[245]^x[235]^x[224]^x[218]^x[217]^x[208]^x[206]^x[197]^x[191]^x[190]^x[181]^x[179]^x[170]^x[130]^x[119]^x[118]^x[117]^x[107]^x[106]^x[103]^x[97]^x[81]^x[75]^x[53]^x[52]^x[51]^x[44]^x[43]^x[33]^x[32];
	y[30]=x[382]^x[381]^x[370]^x[363]^x[362]^x[358]^x[352]^x[350]^x[349]^x[344]^x[343]^x[340]^x[338]^x[334]^x[332]^x[329]^x[323]^x[315]^x[304]^x[286]^x[280]^x[278]^x[277]^x[276]^x[272]^x[271]^x[270]^x[266]^x[265]^x[261]^x[260]^x[259]^x[256]^x[255]^x[254]^x[244]^x[190]^x[189]^x[180]^x[178]^x[169]^x[118]^x[117]^x[116]^x[106]^x[105]^x[102]^x[96]^x[80]^x[74]^x[62]^x[50]^x[43]^x[42]^x[32];
	y[29]=x[383]^x[381]^x[380]^x[369]^x[361]^x[357]^x[349]^x[348]^x[343]^x[342]^x[339]^x[337]^x[333]^x[331]^x[328]^x[322]^x[314]^x[303]^x[287]^x[285]^x[281]^x[279]^x[277]^x[276]^x[275]^x[271]^x[270]^x[269]^x[266]^x[265]^x[264]^x[260]^x[259]^x[258]^x[254]^x[253]^x[243]^x[189]^x[188]^x[179]^x[177]^x[168]^x[139]^x[128]^x[127]^x[117]^x[116]^x[115]^x[106]^x[105]^x[104]^x[101]^x[79]^x[73]^x[63]^x[61]^x[51]^x[49]^x[41];
	y[28]=x[382]^x[380]^x[379]^x[368]^x[360]^x[356]^x[348]^x[347]^x[342]^x[341]^x[338]^x[336]^x[332]^x[330]^x[327]^x[321]^x[313]^x[302]^x[286]^x[284]^x[280]^x[278]^x[276]^x[275]^x[274]^x[270]^x[269]^x[268]^x[265]^x[264]^x[263]^x[259]^x[258]^x[257]^x[253]^x[252]^x[242]^x[188]^x[187]^x[178]^x[176]^x[167]^x[138]^x[126]^x[116]^x[115]^x[114]^x[105]^x[104]^x[103]^x[100]^x[78]^x[72]^x[62]^x[60]^x[50]^x[48]^x[40];
	y[27]=x[381]^x[379]^x[378]^x[367]^x[359]^x[355]^x[347]^x[346]^x[341]^x[340]^x[337]^x[335]^x[331]^x[329]^x[326]^x[320]^x[312]^x[301]^x[285]^x[283]^x[279]^x[277]^x[275]^x[274]^x[273]^x[269]^x[268]^x[267]^x[264]^x[263]^x[262]^x[258]^x[257]^x[256]^x[252]^x[251]^x[241]^x[187]^x[186]^x[177]^x[175]^x[166]^x[137]^x[125]^x[115]^x[114]^x[113]^x[104]^x[103]^x[102]^x[99]^x[77]^x[71]^x[61]^x[59]^x[49]^x[47]^x[39];
	y[26]=x[383]^x[382]^x[380]^x[376]^x[373]^x[372]^x[371]^x[367]^x[365]^x[363]^x[358]^x[354]^x[352]^x[351]^x[346]^x[345]^x[340]^x[339]^x[336]^x[334]^x[328]^x[325]^x[311]^x[300]^x[287]^x[284]^x[282]^x[277]^x[276]^x[274]^x[273]^x[272]^x[268]^x[263]^x[262]^x[261]^x[257]^x[256]^x[251]^x[250]^x[240]^x[223]^x[222]^x[213]^x[212]^x[211]^x[203]^x[192]^x[186]^x[185]^x[176]^x[174]^x[165]^x[157]^x[124]^x[114]^x[113]^x[112]^x[103]^x[102]^x[101]^x[98]^x[76]^x[70]^x[60]^x[48]^x[46]^x[38]^x[37]^x[31]^x[10];
	y[25]=x[381]^x[379]^x[377]^x[376]^x[375]^x[372]^x[370]^x[366]^x[365]^x[364]^x[357]^x[353]^x[350]^x[345]^x[344]^x[339]^x[338]^x[335]^x[333]^x[327]^x[324]^x[310]^x[299]^x[287]^x[286]^x[283]^x[281]^x[277]^x[276]^x[275]^x[273]^x[272]^x[271]^x[267]^x[262]^x[261]^x[260]^x[256]^x[250]^x[249]^x[239]^x[221]^x[212]^x[210]^x[185]^x[184]^x[175]^x[173]^x[164]^x[156]^x[135]^x[123]^x[113]^x[112]^x[111]^x[102]^x[101]^x[100]^x[97]^x[75]^x[69]^x[59]^x[57]^x[47]^x[45]^x[37]^x[30]^x[9];
	y[24]=x[380]^x[378]^x[376]^x[375]^x[374]^x[371]^x[369]^x[365]^x[364]^x[363]^x[356]^x[352]^x[349]^x[344]^x[343]^x[338]^x[337]^x[334]^x[332]^x[326]^x[323]^x[309]^x[298]^x[287]^x[286]^x[285]^x[282]^x[280]^x[276]^x[275]^x[274]^x[272]^x[271]^x[270]^x[261]^x[260]^x[259]^x[249]^x[248]^x[238]^x[220]^x[211]^x[209]^x[184]^x[183]^x[174]^x[172]^x[163]^x[155]^x[134]^x[122]^x[112]^x[111]^x[110]^x[101]^x[100]^x[99]^x[96]^x[74]^x[68]^x[58]^x[56]^x[46]^x[44]^x[36]^x[29]^x[8];
	y[23]=x[379]^x[377]^x[375]^x[373]^x[370]^x[368]^x[364]^x[362]^x[355]^x[348]^x[343]^x[342]^x[337]^x[336]^x[333]^x[331]^x[325]^x[322]^x[308]^x[297]^x[286]^x[285]^x[284]^x[281]^x[279]^x[275]^x[274]^x[273]^x[271]^x[270]^x[269]^x[260]^x[259]^x[258]^x[248]^x[247]^x[237]^x[219]^x[210]^x[208]^x[183]^x[182]^x[173]^x[171]^x[162]^x[154]^x[121]^x[111]^x[110]^x[109]^x[100]^x[99]^x[98]^x[73]^x[67]^x[57]^x[55]^x[45]^x[43]^x[35]^x[28]^x[7];
	y[22]=x[378]^x[376]^x[374]^x[372]^x[369]^x[367]^x[363]^x[361]^x[354]^x[347]^x[342]^x[341]^x[336]^x[335]^x[332]^x[330]^x[324]^x[321]^x[307]^x[296]^x[285]^x[284]^x[283]^x[280]^x[278]^x[274]^x[273]^x[272]^x[270]^x[269]^x[268]^x[259]^x[258]^x[257]^x[247]^x[246]^x[236]^x[218]^x[209]^x[207]^x[182]^x[181]^x[172]^x[170]^x[161]^x[153]^x[120]^x[110]^x[109]^x[108]^x[99]^x[98]^x[97]^x[72]^x[66]^x[56]^x[54]^x[44]^x[42]^x[34]^x[27]^x[6];
	y[21]=x[377]^x[375]^x[373]^x[371]^x[368]^x[366]^x[363]^x[360]^x[353]^x[352]^x[346]^x[341]^x[340]^x[335]^x[334]^x[331]^x[329]^x[323]^x[320]^x[306]^x[295]^x[284]^x[283]^x[282]^x[279]^x[277]^x[273]^x[272]^x[271]^x[269]^x[268]^x[267]^x[258]^x[257]^x[256]^x[246]^x[245]^x[235]^x[217]^x[208]^x[206]^x[181]^x[180]^x[171]^x[169]^x[160]^x[152]^x[119]^x[109]^x[108]^x[107]^x[98]^x[97]^x[96]^x[71]^x[65]^x[55]^x[53]^x[42]^x[41]^x[33]^x[32]^x[26]^x[5];
	y[20]=x[383]^x[382]^x[378]^x[377]^x[374]^x[372]^x[370]^x[366]^x[361]^x[352]^x[351]^x[345]^x[340]^x[339]^x[334]^x[333]^x[328]^x[322]^x[305]^x[294]^x[287]^x[283]^x[282]^x[281]^x[278]^x[276]^x[270]^x[268]^x[267]^x[261]^x[257]^x[256]^x[245]^x[244]^x[234]^x[218]^x[217]^x[206]^x[191]^x[180]^x[179]^x[168]^x[130]^x[127]^x[118]^x[108]^x[107]^x[97]^x[96]^x[70]^x[64]^x[63]^x[62]^x[54]^x[42]^x[41]^x[40]^x[32];
	y[19]=x[383]^x[381]^x[373]^x[370]^x[369]^x[362]^x[360]^x[359]^x[350]^x[344]^x[339]^x[338]^x[333]^x[332]^x[327]^x[321]^x[304]^x[293]^x[287]^x[286]^x[282]^x[281]^x[280]^x[277]^x[275]^x[271]^x[269]^x[267]^x[256]^x[244]^x[243]^x[233]^x[190]^x[179]^x[178]^x[167]^x[127]^x[126]^x[117]^x[107]^x[96]^x[69]^x[63]^x[61]^x[53]^x[51]^x[42]^x[41]^x[40]^x[39];
	y[18]=x[382]^x[380]^x[372]^x[369]^x[368]^x[361]^x[359]^x[358]^x[349]^x[343]^x[338]^x[337]^x[332]^x[331]^x[326]^x[320]^x[303]^x[292]^x[287]^x[286]^x[285]^x[281]^x[280]^x[279]^x[276]^x[274]^x[270]^x[268]^x[243]^x[242]^x[232]^x[189]^x[178]^x[177]^x[166]^x[127]^x[126]^x[125]^x[116]^x[68]^x[62]^x[60]^x[52]^x[50]^x[41]^x[40]^x[39]^x[38];
	y[17]=x[381]^x[379]^x[374]^x[373]^x[371]^x[362]^x[360]^x[358]^x[356]^x[352]^x[348]^x[342]^x[337]^x[336]^x[331]^x[325]^x[302]^x[291]^x[286]^x[285]^x[284]^x[280]^x[279]^x[278]^x[275]^x[273]^x[269]^x[267]^x[242]^x[241]^x[231]^x[214]^x[213]^x[202]^x[192]^x[188]^x[177]^x[176]^x[165]^x[126]^x[125]^x[124]^x[115]^x[67]^x[61]^x[59]^x[51]^x[49]^x[40]^x[39]^x[38]^x[37];
	y[16]=x[380]^x[378]^x[372]^x[370]^x[367]^x[361]^x[359]^x[357]^x[356]^x[355]^x[347]^x[341]^x[336]^x[335]^x[330]^x[324]^x[301]^x[290]^x[285]^x[284]^x[283]^x[279]^x[278]^x[277]^x[274]^x[272]^x[268]^x[266]^x[241]^x[240]^x[230]^x[212]^x[201]^x[187]^x[176]^x[175]^x[164]^x[125]^x[124]^x[123]^x[114]^x[66]^x[60]^x[58]^x[50]^x[48]^x[39]^x[38]^x[37]^x[36];
	y[15]=x[379]^x[377]^x[373]^x[371]^x[369]^x[367]^x[366]^x[362]^x[360]^x[358]^x[355]^x[354]^x[346]^x[340]^x[335]^x[334]^x[329]^x[323]^x[300]^x[289]^x[284]^x[283]^x[282]^x[278]^x[277]^x[276]^x[273]^x[271]^x[266]^x[265]^x[256]^x[240]^x[239]^x[229]^x[213]^x[211]^x[202]^x[200]^x[186]^x[175]^x[174]^x[163]^x[124]^x[123]^x[122]^x[113]^x[65]^x[59]^x[57]^x[49]^x[47]^x[38]^x[37]^x[36]^x[35];
	y[14]=x[378]^x[376]^x[372]^x[370]^x[368]^x[366]^x[365]^x[361]^x[359]^x[357]^x[354]^x[353]^x[345]^x[339]^x[334]^x[333]^x[328]^x[322]^x[299]^x[288]^x[283]^x[282]^x[281]^x[277]^x[276]^x[275]^x[272]^x[270]^x[266]^x[265]^x[264]^x[239]^x[238]^x[228]^x[212]^x[210]^x[201]^x[199]^x[185]^x[174]^x[173]^x[162]^x[123]^x[122]^x[121]^x[112]^x[64]^x[58]^x[56]^x[48]^x[46]^x[37]^x[36]^x[35]^x[34];
	y[13]=x[377]^x[375]^x[371]^x[369]^x[367]^x[365]^x[364]^x[360]^x[358]^x[356]^x[353]^x[352]^x[344]^x[338]^x[333]^x[332]^x[327]^x[321]^x[282]^x[281]^x[280]^x[276]^x[275]^x[274]^x[271]^x[269]^x[265]^x[264]^x[263]^x[238]^x[237]^x[227]^x[211]^x[209]^x[200]^x[198]^x[184]^x[173]^x[172]^x[161]^x[122]^x[121]^x[120]^x[111]^x[57]^x[55]^x[47]^x[45]^x[36]^x[35]^x[34]^x[33];
	y[12]=x[376]^x[374]^x[370]^x[368]^x[366]^x[364]^x[359]^x[357]^x[355]^x[343]^x[337]^x[332]^x[331]^x[326]^x[320]^x[281]^x[280]^x[279]^x[275]^x[274]^x[273]^x[270]^x[268]^x[264]^x[263]^x[262]^x[237]^x[236]^x[226]^x[210]^x[208]^x[199]^x[197]^x[183]^x[172]^x[171]^x[160]^x[121]^x[120]^x[119]^x[110]^x[56]^x[54]^x[46]^x[44]^x[35]^x[34]^x[33]^x[32];
	y[11]=x[375]^x[374]^x[369]^x[368]^x[365]^x[358]^x[357]^x[354]^x[342]^x[336]^x[331]^x[325]^x[280]^x[279]^x[278]^x[274]^x[273]^x[272]^x[269]^x[267]^x[263]^x[262]^x[261]^x[236]^x[235]^x[225]^x[209]^x[208]^x[198]^x[197]^x[182]^x[171]^x[120]^x[119]^x[118]^x[109]^x[55]^x[54]^x[45]^x[34]^x[33]^x[32];
	y[10]=x[374]^x[368]^x[364]^x[362]^x[357]^x[353]^x[341]^x[335]^x[330]^x[324]^x[279]^x[278]^x[277]^x[273]^x[272]^x[271]^x[268]^x[266]^x[262]^x[261]^x[260]^x[235]^x[234]^x[224]^x[208]^x[197]^x[181]^x[170]^x[119]^x[118]^x[117]^x[108]^x[54]^x[44]^x[42]^x[33]^x[32];
	y[9]=x[381]^x[373]^x[372]^x[371]^x[363]^x[359]^x[352]^x[340]^x[334]^x[329]^x[323]^x[282]^x[278]^x[277]^x[276]^x[272]^x[271]^x[270]^x[267]^x[265]^x[261]^x[259]^x[255]^x[233]^x[180]^x[169]^x[118]^x[117]^x[116]^x[107]^x[53]^x[52]^x[51]^x[43]^x[41]^x[32];
	y[8]=x[383]^x[380]^x[372]^x[371]^x[370]^x[358]^x[339]^x[333]^x[328]^x[322]^x[277]^x[276]^x[275]^x[271]^x[270]^x[269]^x[266]^x[264]^x[260]^x[258]^x[254]^x[232]^x[179]^x[168]^x[117]^x[116]^x[115]^x[106]^x[63]^x[52]^x[50]^x[40];
	y[7]=x[382]^x[379]^x[371]^x[370]^x[369]^x[357]^x[338]^x[332]^x[327]^x[321]^x[276]^x[275]^x[274]^x[270]^x[269]^x[268]^x[265]^x[263]^x[259]^x[257]^x[253]^x[231]^x[178]^x[167]^x[138]^x[116]^x[115]^x[114]^x[105]^x[62]^x[51]^x[49]^x[39];
	y[6]=x[381]^x[378]^x[370]^x[369]^x[368]^x[356]^x[337]^x[331]^x[326]^x[320]^x[275]^x[274]^x[273]^x[269]^x[268]^x[267]^x[264]^x[262]^x[258]^x[256]^x[252]^x[230]^x[177]^x[166]^x[137]^x[115]^x[114]^x[113]^x[104]^x[61]^x[50]^x[48]^x[38];
	y[5]=x[380]^x[377]^x[374]^x[369]^x[367]^x[357]^x[355]^x[352]^x[336]^x[325]^x[278]^x[274]^x[273]^x[272]^x[263]^x[261]^x[256]^x[251]^x[229]^x[214]^x[192]^x[176]^x[165]^x[136]^x[114]^x[113]^x[112]^x[103]^x[60]^x[49]^x[47]^x[10];
	y[4]=x[379]^x[376]^x[373]^x[368]^x[366]^x[362]^x[356]^x[354]^x[335]^x[324]^x[273]^x[272]^x[271]^x[262]^x[260]^x[250]^x[228]^x[213]^x[202]^x[175]^x[164]^x[135]^x[113]^x[112]^x[111]^x[102]^x[59]^x[48]^x[46]^x[36]^x[9];
	y[3]=x[378]^x[375]^x[372]^x[367]^x[365]^x[361]^x[355]^x[353]^x[334]^x[323]^x[272]^x[271]^x[270]^x[261]^x[259]^x[249]^x[227]^x[212]^x[201]^x[174]^x[163]^x[134]^x[112]^x[111]^x[110]^x[101]^x[58]^x[47]^x[45]^x[35]^x[8];
	y[2]=x[377]^x[374]^x[371]^x[366]^x[364]^x[360]^x[354]^x[352]^x[333]^x[322]^x[271]^x[270]^x[269]^x[260]^x[258]^x[248]^x[226]^x[211]^x[200]^x[173]^x[162]^x[133]^x[111]^x[110]^x[109]^x[100]^x[57]^x[46]^x[44]^x[34]^x[7];
	y[1]=x[376]^x[370]^x[365]^x[363]^x[359]^x[353]^x[332]^x[321]^x[270]^x[269]^x[268]^x[259]^x[257]^x[247]^x[225]^x[210]^x[199]^x[172]^x[161]^x[110]^x[109]^x[108]^x[99]^x[56]^x[45]^x[43]^x[33]^x[6];
	y[0]=x[375]^x[369]^x[364]^x[363]^x[358]^x[331]^x[320]^x[269]^x[268]^x[267]^x[258]^x[256]^x[246]^x[224]^x[209]^x[198]^x[171]^x[160]^x[109]^x[108]^x[107]^x[98]^x[55]^x[44]^x[43]^x[5];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint57(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[346]^x[345]^x[341]^x[336]^x[334]^x[332]^x[331]^x[330]^x[327]^x[325]^x[321]^x[319]^x[318]^x[313]^x[312]^x[309]^x[307]^x[303]^x[301]^x[298]^x[292]^x[284]^x[273]^x[255]^x[251]^x[250]^x[249]^x[247]^x[246]^x[245]^x[241]^x[239]^x[235]^x[234]^x[230]^x[229]^x[228]^x[225]^x[223]^x[213]^x[203]^x[192]^x[186]^x[185]^x[176]^x[174]^x[165]^x[159]^x[158]^x[149]^x[147]^x[138]^x[98]^x[87]^x[86]^x[85]^x[75]^x[74]^x[71]^x[65]^x[49]^x[43]^x[21]^x[20]^x[19]^x[12]^x[11]^x[1]^x[0];
	y[30]=x[350]^x[349]^x[338]^x[331]^x[330]^x[326]^x[320]^x[318]^x[317]^x[312]^x[311]^x[308]^x[306]^x[302]^x[300]^x[297]^x[291]^x[283]^x[272]^x[254]^x[248]^x[246]^x[245]^x[244]^x[240]^x[239]^x[238]^x[234]^x[233]^x[229]^x[228]^x[227]^x[224]^x[223]^x[222]^x[212]^x[158]^x[157]^x[148]^x[146]^x[137]^x[86]^x[85]^x[84]^x[74]^x[73]^x[70]^x[64]^x[48]^x[42]^x[30]^x[18]^x[11]^x[10]^x[0];
	y[29]=x[351]^x[349]^x[348]^x[337]^x[329]^x[325]^x[317]^x[316]^x[311]^x[310]^x[307]^x[305]^x[301]^x[299]^x[296]^x[290]^x[282]^x[271]^x[255]^x[253]^x[249]^x[247]^x[245]^x[244]^x[243]^x[239]^x[238]^x[237]^x[234]^x[233]^x[232]^x[228]^x[227]^x[226]^x[222]^x[221]^x[211]^x[157]^x[156]^x[147]^x[145]^x[136]^x[107]^x[96]^x[95]^x[85]^x[84]^x[83]^x[74]^x[73]^x[72]^x[69]^x[47]^x[41]^x[31]^x[29]^x[19]^x[17]^x[9];
	y[28]=x[350]^x[348]^x[347]^x[336]^x[328]^x[324]^x[316]^x[315]^x[310]^x[309]^x[306]^x[304]^x[300]^x[298]^x[295]^x[289]^x[281]^x[270]^x[254]^x[252]^x[248]^x[246]^x[244]^x[243]^x[242]^x[238]^x[237]^x[236]^x[233]^x[232]^x[231]^x[227]^x[226]^x[225]^x[221]^x[220]^x[210]^x[156]^x[155]^x[146]^x[144]^x[135]^x[106]^x[94]^x[84]^x[83]^x[82]^x[73]^x[72]^x[71]^x[68]^x[46]^x[40]^x[30]^x[28]^x[18]^x[16]^x[8];
	y[27]=x[349]^x[347]^x[346]^x[335]^x[327]^x[323]^x[315]^x[314]^x[309]^x[308]^x[305]^x[303]^x[299]^x[297]^x[294]^x[288]^x[280]^x[269]^x[253]^x[251]^x[247]^x[245]^x[243]^x[242]^x[241]^x[237]^x[236]^x[235]^x[232]^x[231]^x[230]^x[226]^x[225]^x[224]^x[220]^x[219]^x[209]^x[155]^x[154]^x[145]^x[143]^x[134]^x[105]^x[93]^x[83]^x[82]^x[81]^x[72]^x[71]^x[70]^x[67]^x[45]^x[39]^x[29]^x[27]^x[17]^x[15]^x[7];
	y[26]=x[383]^x[351]^x[350]^x[348]^x[344]^x[341]^x[340]^x[339]^x[335]^x[333]^x[331]^x[326]^x[322]^x[320]^x[319]^x[314]^x[313]^x[308]^x[307]^x[304]^x[302]^x[296]^x[293]^x[279]^x[268]^x[255]^x[252]^x[250]^x[245]^x[244]^x[242]^x[241]^x[240]^x[236]^x[231]^x[230]^x[229]^x[225]^x[224]^x[219]^x[218]^x[208]^x[191]^x[190]^x[181]^x[180]^x[179]^x[171]^x[160]^x[159]^x[154]^x[144]^x[142]^x[138]^x[133]^x[132]^x[125]^x[92]^x[82]^x[81]^x[80]^x[71]^x[70]^x[69]^x[66]^x[44]^x[38]^x[28]^x[16]^x[14]^x[6]^x[5];
	y[25]=x[382]^x[349]^x[347]^x[345]^x[344]^x[343]^x[340]^x[338]^x[334]^x[333]^x[332]^x[325]^x[321]^x[318]^x[313]^x[312]^x[307]^x[306]^x[303]^x[301]^x[295]^x[292]^x[278]^x[267]^x[255]^x[254]^x[251]^x[249]^x[245]^x[244]^x[243]^x[241]^x[240]^x[239]^x[235]^x[230]^x[229]^x[228]^x[224]^x[218]^x[217]^x[207]^x[189]^x[180]^x[178]^x[158]^x[153]^x[143]^x[141]^x[137]^x[132]^x[131]^x[124]^x[103]^x[91]^x[81]^x[80]^x[79]^x[70]^x[69]^x[68]^x[65]^x[43]^x[37]^x[27]^x[25]^x[15]^x[13]^x[5];
	y[24]=x[381]^x[348]^x[346]^x[344]^x[343]^x[342]^x[339]^x[337]^x[333]^x[332]^x[331]^x[324]^x[320]^x[317]^x[312]^x[311]^x[306]^x[305]^x[302]^x[300]^x[294]^x[291]^x[277]^x[266]^x[255]^x[254]^x[253]^x[250]^x[248]^x[244]^x[243]^x[242]^x[240]^x[239]^x[238]^x[229]^x[228]^x[227]^x[217]^x[216]^x[206]^x[188]^x[179]^x[177]^x[157]^x[152]^x[142]^x[140]^x[136]^x[131]^x[130]^x[123]^x[102]^x[90]^x[80]^x[79]^x[78]^x[69]^x[68]^x[67]^x[64]^x[42]^x[36]^x[26]^x[24]^x[14]^x[12]^x[4];
	y[23]=x[380]^x[347]^x[345]^x[343]^x[341]^x[338]^x[336]^x[332]^x[330]^x[323]^x[316]^x[311]^x[310]^x[305]^x[304]^x[301]^x[299]^x[293]^x[290]^x[276]^x[265]^x[254]^x[253]^x[252]^x[249]^x[247]^x[243]^x[242]^x[241]^x[239]^x[238]^x[237]^x[228]^x[227]^x[226]^x[216]^x[215]^x[205]^x[187]^x[178]^x[176]^x[156]^x[151]^x[141]^x[139]^x[135]^x[130]^x[129]^x[122]^x[89]^x[79]^x[78]^x[77]^x[68]^x[67]^x[66]^x[41]^x[35]^x[25]^x[23]^x[13]^x[11]^x[3];
	y[22]=x[379]^x[346]^x[344]^x[342]^x[340]^x[337]^x[335]^x[331]^x[329]^x[322]^x[315]^x[310]^x[309]^x[304]^x[303]^x[300]^x[298]^x[292]^x[289]^x[275]^x[264]^x[253]^x[252]^x[251]^x[248]^x[246]^x[242]^x[241]^x[240]^x[238]^x[237]^x[236]^x[227]^x[226]^x[225]^x[215]^x[214]^x[204]^x[186]^x[177]^x[175]^x[155]^x[150]^x[140]^x[138]^x[134]^x[129]^x[128]^x[121]^x[88]^x[78]^x[77]^x[76]^x[67]^x[66]^x[65]^x[40]^x[34]^x[24]^x[22]^x[12]^x[10]^x[2];
	y[21]=x[378]^x[345]^x[343]^x[341]^x[339]^x[336]^x[334]^x[331]^x[328]^x[321]^x[320]^x[314]^x[309]^x[308]^x[303]^x[302]^x[299]^x[297]^x[291]^x[288]^x[274]^x[263]^x[252]^x[251]^x[250]^x[247]^x[245]^x[241]^x[240]^x[239]^x[237]^x[236]^x[235]^x[226]^x[225]^x[224]^x[214]^x[213]^x[203]^x[185]^x[176]^x[174]^x[154]^x[149]^x[139]^x[137]^x[133]^x[128]^x[120]^x[87]^x[77]^x[76]^x[75]^x[66]^x[65]^x[64]^x[39]^x[33]^x[23]^x[21]^x[10]^x[9]^x[1]^x[0];
	y[20]=x[351]^x[350]^x[346]^x[345]^x[342]^x[340]^x[338]^x[334]^x[329]^x[320]^x[319]^x[313]^x[308]^x[307]^x[302]^x[301]^x[296]^x[290]^x[273]^x[262]^x[255]^x[251]^x[250]^x[249]^x[246]^x[244]^x[238]^x[236]^x[235]^x[229]^x[225]^x[224]^x[213]^x[212]^x[202]^x[186]^x[185]^x[174]^x[159]^x[148]^x[147]^x[136]^x[98]^x[95]^x[86]^x[76]^x[75]^x[65]^x[64]^x[38]^x[32]^x[31]^x[30]^x[22]^x[10]^x[9]^x[8]^x[0];
	y[19]=x[351]^x[349]^x[341]^x[338]^x[337]^x[330]^x[328]^x[327]^x[318]^x[312]^x[307]^x[306]^x[301]^x[300]^x[295]^x[289]^x[272]^x[261]^x[255]^x[254]^x[250]^x[249]^x[248]^x[245]^x[243]^x[239]^x[237]^x[235]^x[224]^x[212]^x[211]^x[201]^x[158]^x[147]^x[146]^x[135]^x[95]^x[94]^x[85]^x[75]^x[64]^x[37]^x[31]^x[29]^x[21]^x[19]^x[10]^x[9]^x[8]^x[7];
	y[18]=x[350]^x[348]^x[340]^x[337]^x[336]^x[329]^x[327]^x[326]^x[317]^x[311]^x[306]^x[305]^x[300]^x[299]^x[294]^x[288]^x[271]^x[260]^x[255]^x[254]^x[253]^x[249]^x[248]^x[247]^x[244]^x[242]^x[238]^x[236]^x[211]^x[210]^x[200]^x[157]^x[146]^x[145]^x[134]^x[95]^x[94]^x[93]^x[84]^x[36]^x[30]^x[28]^x[20]^x[18]^x[9]^x[8]^x[7]^x[6];
	y[17]=x[349]^x[347]^x[342]^x[341]^x[339]^x[330]^x[328]^x[326]^x[324]^x[320]^x[316]^x[310]^x[305]^x[304]^x[299]^x[293]^x[270]^x[259]^x[254]^x[253]^x[252]^x[248]^x[247]^x[246]^x[243]^x[241]^x[237]^x[235]^x[210]^x[209]^x[199]^x[182]^x[181]^x[170]^x[160]^x[156]^x[145]^x[144]^x[133]^x[94]^x[93]^x[92]^x[83]^x[35]^x[29]^x[27]^x[19]^x[17]^x[8]^x[7]^x[6]^x[5];
	y[16]=x[348]^x[346]^x[340]^x[338]^x[335]^x[329]^x[327]^x[325]^x[324]^x[323]^x[315]^x[309]^x[304]^x[303]^x[298]^x[292]^x[269]^x[258]^x[253]^x[252]^x[251]^x[247]^x[246]^x[245]^x[242]^x[240]^x[236]^x[234]^x[209]^x[208]^x[198]^x[180]^x[169]^x[155]^x[144]^x[143]^x[132]^x[93]^x[92]^x[91]^x[82]^x[34]^x[28]^x[26]^x[18]^x[16]^x[7]^x[6]^x[5]^x[4];
	y[15]=x[347]^x[345]^x[341]^x[339]^x[337]^x[335]^x[334]^x[330]^x[328]^x[326]^x[323]^x[322]^x[314]^x[308]^x[303]^x[302]^x[297]^x[291]^x[268]^x[257]^x[252]^x[251]^x[250]^x[246]^x[245]^x[244]^x[241]^x[239]^x[234]^x[233]^x[224]^x[208]^x[207]^x[197]^x[181]^x[179]^x[170]^x[168]^x[154]^x[143]^x[142]^x[131]^x[92]^x[91]^x[90]^x[81]^x[33]^x[27]^x[25]^x[17]^x[15]^x[6]^x[5]^x[4]^x[3];
	y[14]=x[346]^x[344]^x[340]^x[338]^x[336]^x[334]^x[333]^x[329]^x[327]^x[325]^x[322]^x[321]^x[313]^x[307]^x[302]^x[301]^x[296]^x[290]^x[267]^x[256]^x[251]^x[250]^x[249]^x[245]^x[244]^x[243]^x[240]^x[238]^x[234]^x[233]^x[232]^x[207]^x[206]^x[196]^x[180]^x[178]^x[169]^x[167]^x[153]^x[142]^x[141]^x[130]^x[91]^x[90]^x[89]^x[80]^x[32]^x[26]^x[24]^x[16]^x[14]^x[5]^x[4]^x[3]^x[2];
	y[13]=x[345]^x[343]^x[339]^x[337]^x[335]^x[333]^x[332]^x[328]^x[326]^x[324]^x[321]^x[320]^x[312]^x[306]^x[301]^x[300]^x[295]^x[289]^x[250]^x[249]^x[248]^x[244]^x[243]^x[242]^x[239]^x[237]^x[233]^x[232]^x[231]^x[206]^x[205]^x[195]^x[179]^x[177]^x[168]^x[166]^x[152]^x[141]^x[140]^x[129]^x[90]^x[89]^x[88]^x[79]^x[25]^x[23]^x[15]^x[13]^x[4]^x[3]^x[2]^x[1];
	y[12]=x[344]^x[342]^x[338]^x[336]^x[334]^x[332]^x[327]^x[325]^x[323]^x[311]^x[305]^x[300]^x[299]^x[294]^x[288]^x[249]^x[248]^x[247]^x[243]^x[242]^x[241]^x[238]^x[236]^x[232]^x[231]^x[230]^x[205]^x[204]^x[194]^x[178]^x[176]^x[167]^x[165]^x[151]^x[140]^x[139]^x[128]^x[89]^x[88]^x[87]^x[78]^x[24]^x[22]^x[14]^x[12]^x[3]^x[2]^x[1]^x[0];
	y[11]=x[343]^x[342]^x[337]^x[336]^x[333]^x[326]^x[325]^x[322]^x[310]^x[304]^x[299]^x[293]^x[248]^x[247]^x[246]^x[242]^x[241]^x[240]^x[237]^x[235]^x[231]^x[230]^x[229]^x[204]^x[203]^x[193]^x[177]^x[176]^x[166]^x[165]^x[150]^x[139]^x[88]^x[87]^x[86]^x[77]^x[23]^x[22]^x[13]^x[2]^x[1]^x[0];
	y[10]=x[342]^x[336]^x[332]^x[330]^x[325]^x[321]^x[309]^x[303]^x[298]^x[292]^x[247]^x[246]^x[245]^x[241]^x[240]^x[239]^x[236]^x[234]^x[230]^x[229]^x[228]^x[203]^x[202]^x[192]^x[176]^x[165]^x[149]^x[138]^x[87]^x[86]^x[85]^x[76]^x[22]^x[12]^x[10]^x[1]^x[0];
	y[9]=x[349]^x[341]^x[340]^x[339]^x[331]^x[327]^x[320]^x[308]^x[302]^x[297]^x[291]^x[250]^x[246]^x[245]^x[244]^x[240]^x[239]^x[238]^x[235]^x[233]^x[229]^x[227]^x[223]^x[201]^x[148]^x[137]^x[86]^x[85]^x[84]^x[75]^x[21]^x[20]^x[19]^x[11]^x[9]^x[0];
	y[8]=x[351]^x[348]^x[340]^x[339]^x[338]^x[326]^x[307]^x[301]^x[296]^x[290]^x[245]^x[244]^x[243]^x[239]^x[238]^x[237]^x[234]^x[232]^x[228]^x[226]^x[222]^x[200]^x[147]^x[136]^x[85]^x[84]^x[83]^x[74]^x[31]^x[20]^x[18]^x[8];
	y[7]=x[350]^x[347]^x[339]^x[338]^x[337]^x[325]^x[306]^x[300]^x[295]^x[289]^x[244]^x[243]^x[242]^x[238]^x[237]^x[236]^x[233]^x[231]^x[227]^x[225]^x[221]^x[199]^x[146]^x[135]^x[106]^x[84]^x[83]^x[82]^x[73]^x[30]^x[19]^x[17]^x[7];
	y[6]=x[349]^x[346]^x[338]^x[337]^x[336]^x[324]^x[305]^x[299]^x[294]^x[288]^x[243]^x[242]^x[241]^x[237]^x[236]^x[235]^x[232]^x[230]^x[226]^x[224]^x[220]^x[198]^x[145]^x[134]^x[105]^x[83]^x[82]^x[81]^x[72]^x[29]^x[18]^x[16]^x[6];
	y[5]=x[373]^x[362]^x[348]^x[345]^x[342]^x[337]^x[335]^x[325]^x[323]^x[320]^x[304]^x[293]^x[246]^x[242]^x[241]^x[240]^x[231]^x[229]^x[224]^x[219]^x[197]^x[182]^x[160]^x[144]^x[138]^x[133]^x[132]^x[104]^x[82]^x[81]^x[80]^x[71]^x[28]^x[17]^x[15];
	y[4]=x[372]^x[361]^x[347]^x[344]^x[341]^x[336]^x[334]^x[330]^x[324]^x[322]^x[303]^x[292]^x[241]^x[240]^x[239]^x[230]^x[228]^x[218]^x[196]^x[181]^x[170]^x[143]^x[137]^x[132]^x[131]^x[103]^x[81]^x[80]^x[79]^x[70]^x[27]^x[16]^x[14]^x[4];
	y[3]=x[371]^x[360]^x[346]^x[343]^x[340]^x[335]^x[333]^x[329]^x[323]^x[321]^x[302]^x[291]^x[240]^x[239]^x[238]^x[229]^x[227]^x[217]^x[195]^x[180]^x[169]^x[142]^x[136]^x[131]^x[130]^x[102]^x[80]^x[79]^x[78]^x[69]^x[26]^x[15]^x[13]^x[3];
	y[2]=x[370]^x[359]^x[345]^x[342]^x[339]^x[334]^x[332]^x[328]^x[322]^x[320]^x[301]^x[290]^x[239]^x[238]^x[237]^x[228]^x[226]^x[216]^x[194]^x[179]^x[168]^x[141]^x[135]^x[130]^x[129]^x[101]^x[79]^x[78]^x[77]^x[68]^x[25]^x[14]^x[12]^x[2];
	y[1]=x[369]^x[358]^x[344]^x[338]^x[333]^x[331]^x[327]^x[321]^x[300]^x[289]^x[238]^x[237]^x[236]^x[227]^x[225]^x[215]^x[193]^x[178]^x[167]^x[140]^x[134]^x[129]^x[128]^x[78]^x[77]^x[76]^x[67]^x[24]^x[13]^x[11]^x[1];
	y[0]=x[368]^x[357]^x[343]^x[337]^x[332]^x[331]^x[326]^x[299]^x[288]^x[237]^x[236]^x[235]^x[226]^x[224]^x[214]^x[192]^x[177]^x[166]^x[139]^x[133]^x[128]^x[77]^x[76]^x[75]^x[66]^x[23]^x[12]^x[11];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint58(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[375]^x[374]^x[373]^x[372]^x[371]^x[363]^x[353]^x[314]^x[313]^x[309]^x[304]^x[302]^x[300]^x[299]^x[298]^x[295]^x[293]^x[289]^x[287]^x[286]^x[281]^x[280]^x[277]^x[275]^x[271]^x[269]^x[266]^x[260]^x[252]^x[241]^x[223]^x[219]^x[218]^x[217]^x[215]^x[214]^x[213]^x[209]^x[207]^x[203]^x[202]^x[198]^x[197]^x[196]^x[193]^x[191]^x[181]^x[171]^x[160]^x[154]^x[153]^x[149]^x[148]^x[147]^x[144]^x[143]^x[141]^x[140]^x[139]^x[134]^x[129]^x[128]^x[127]^x[126]^x[117]^x[115]^x[106]^x[66]^x[55]^x[54]^x[53]^x[43]^x[42]^x[39]^x[33]^x[17]^x[11];
	y[30]=x[382]^x[381]^x[374]^x[373]^x[372]^x[370]^x[362]^x[361]^x[352]^x[318]^x[317]^x[306]^x[299]^x[298]^x[294]^x[288]^x[286]^x[285]^x[280]^x[279]^x[276]^x[274]^x[270]^x[268]^x[265]^x[259]^x[251]^x[240]^x[222]^x[216]^x[214]^x[213]^x[212]^x[208]^x[207]^x[206]^x[202]^x[201]^x[197]^x[196]^x[195]^x[192]^x[191]^x[190]^x[180]^x[158]^x[152]^x[146]^x[140]^x[139]^x[138]^x[133]^x[132]^x[128]^x[126]^x[125]^x[116]^x[114]^x[105]^x[54]^x[53]^x[52]^x[42]^x[41]^x[38]^x[32]^x[16]^x[10];
	y[29]=x[383]^x[382]^x[381]^x[380]^x[373]^x[372]^x[369]^x[362]^x[361]^x[360]^x[319]^x[317]^x[316]^x[305]^x[297]^x[293]^x[285]^x[284]^x[279]^x[278]^x[275]^x[273]^x[269]^x[267]^x[264]^x[258]^x[250]^x[239]^x[223]^x[221]^x[217]^x[215]^x[213]^x[212]^x[211]^x[207]^x[206]^x[205]^x[202]^x[201]^x[200]^x[196]^x[195]^x[194]^x[190]^x[189]^x[179]^x[159]^x[157]^x[153]^x[151]^x[147]^x[145]^x[141]^x[139]^x[137]^x[131]^x[125]^x[124]^x[115]^x[113]^x[104]^x[75]^x[64]^x[63]^x[53]^x[52]^x[51]^x[42]^x[41]^x[40]^x[37]^x[15]^x[9];
	y[28]=x[382]^x[381]^x[380]^x[379]^x[372]^x[371]^x[368]^x[361]^x[360]^x[359]^x[318]^x[316]^x[315]^x[304]^x[296]^x[292]^x[284]^x[283]^x[278]^x[277]^x[274]^x[272]^x[268]^x[266]^x[263]^x[257]^x[249]^x[238]^x[222]^x[220]^x[216]^x[214]^x[212]^x[211]^x[210]^x[206]^x[205]^x[204]^x[201]^x[200]^x[199]^x[195]^x[194]^x[193]^x[189]^x[188]^x[178]^x[158]^x[156]^x[152]^x[150]^x[146]^x[144]^x[140]^x[138]^x[136]^x[130]^x[124]^x[123]^x[114]^x[112]^x[103]^x[74]^x[62]^x[52]^x[51]^x[50]^x[41]^x[40]^x[39]^x[36]^x[14]^x[8];
	y[27]=x[381]^x[380]^x[379]^x[378]^x[371]^x[370]^x[367]^x[360]^x[359]^x[358]^x[317]^x[315]^x[314]^x[303]^x[295]^x[291]^x[283]^x[282]^x[277]^x[276]^x[273]^x[271]^x[267]^x[265]^x[262]^x[256]^x[248]^x[237]^x[221]^x[219]^x[215]^x[213]^x[211]^x[210]^x[209]^x[205]^x[204]^x[203]^x[200]^x[199]^x[198]^x[194]^x[193]^x[192]^x[188]^x[187]^x[177]^x[157]^x[155]^x[151]^x[149]^x[145]^x[143]^x[139]^x[137]^x[135]^x[129]^x[123]^x[122]^x[113]^x[111]^x[102]^x[73]^x[61]^x[51]^x[50]^x[49]^x[40]^x[39]^x[38]^x[35]^x[13]^x[7];
	y[26]=x[380]^x[379]^x[377]^x[370]^x[369]^x[366]^x[359]^x[358]^x[357]^x[351]^x[319]^x[318]^x[316]^x[312]^x[309]^x[308]^x[307]^x[303]^x[301]^x[299]^x[294]^x[290]^x[288]^x[287]^x[282]^x[281]^x[276]^x[275]^x[272]^x[270]^x[264]^x[261]^x[247]^x[236]^x[223]^x[220]^x[218]^x[213]^x[212]^x[210]^x[209]^x[208]^x[204]^x[199]^x[198]^x[197]^x[193]^x[192]^x[187]^x[186]^x[176]^x[159]^x[158]^x[156]^x[150]^x[149]^x[148]^x[147]^x[144]^x[142]^x[139]^x[138]^x[136]^x[134]^x[133]^x[127]^x[122]^x[112]^x[110]^x[106]^x[101]^x[100]^x[93]^x[60]^x[50]^x[49]^x[48]^x[39]^x[38]^x[37]^x[34]^x[12]^x[6];
	y[25]=x[379]^x[378]^x[377]^x[376]^x[369]^x[368]^x[365]^x[358]^x[357]^x[356]^x[350]^x[317]^x[315]^x[313]^x[312]^x[311]^x[308]^x[306]^x[302]^x[301]^x[300]^x[293]^x[289]^x[286]^x[281]^x[280]^x[275]^x[274]^x[271]^x[269]^x[263]^x[260]^x[246]^x[235]^x[223]^x[222]^x[219]^x[217]^x[213]^x[212]^x[211]^x[209]^x[208]^x[207]^x[203]^x[198]^x[197]^x[196]^x[192]^x[186]^x[185]^x[175]^x[157]^x[155]^x[153]^x[149]^x[148]^x[147]^x[146]^x[143]^x[141]^x[137]^x[135]^x[133]^x[126]^x[121]^x[111]^x[109]^x[105]^x[100]^x[99]^x[92]^x[71]^x[59]^x[49]^x[48]^x[47]^x[38]^x[37]^x[36]^x[33]^x[11]^x[5];
	y[24]=x[378]^x[377]^x[376]^x[375]^x[368]^x[367]^x[364]^x[357]^x[356]^x[355]^x[349]^x[316]^x[314]^x[312]^x[311]^x[310]^x[307]^x[305]^x[301]^x[300]^x[299]^x[292]^x[288]^x[285]^x[280]^x[279]^x[274]^x[273]^x[270]^x[268]^x[262]^x[259]^x[245]^x[234]^x[223]^x[222]^x[221]^x[218]^x[216]^x[212]^x[211]^x[210]^x[208]^x[207]^x[206]^x[197]^x[196]^x[195]^x[185]^x[184]^x[174]^x[156]^x[154]^x[152]^x[148]^x[147]^x[146]^x[145]^x[142]^x[140]^x[136]^x[134]^x[132]^x[125]^x[120]^x[110]^x[108]^x[104]^x[99]^x[98]^x[91]^x[70]^x[58]^x[48]^x[47]^x[46]^x[37]^x[36]^x[35]^x[32]^x[10]^x[4];
	y[23]=x[377]^x[376]^x[375]^x[374]^x[367]^x[366]^x[363]^x[356]^x[355]^x[354]^x[348]^x[315]^x[313]^x[311]^x[309]^x[306]^x[304]^x[300]^x[298]^x[291]^x[284]^x[279]^x[278]^x[273]^x[272]^x[269]^x[267]^x[261]^x[258]^x[244]^x[233]^x[222]^x[221]^x[220]^x[217]^x[215]^x[211]^x[210]^x[209]^x[207]^x[206]^x[205]^x[196]^x[195]^x[194]^x[184]^x[183]^x[173]^x[155]^x[153]^x[151]^x[147]^x[146]^x[145]^x[144]^x[141]^x[139]^x[135]^x[133]^x[131]^x[124]^x[119]^x[109]^x[107]^x[103]^x[98]^x[97]^x[90]^x[57]^x[47]^x[46]^x[45]^x[36]^x[35]^x[34]^x[9]^x[3];
	y[22]=x[376]^x[375]^x[374]^x[373]^x[366]^x[365]^x[362]^x[355]^x[354]^x[353]^x[347]^x[314]^x[312]^x[310]^x[308]^x[305]^x[303]^x[299]^x[297]^x[290]^x[283]^x[278]^x[277]^x[272]^x[271]^x[268]^x[266]^x[260]^x[257]^x[243]^x[232]^x[221]^x[220]^x[219]^x[216]^x[214]^x[210]^x[209]^x[208]^x[206]^x[205]^x[204]^x[195]^x[194]^x[193]^x[183]^x[182]^x[172]^x[154]^x[152]^x[150]^x[146]^x[145]^x[144]^x[143]^x[140]^x[138]^x[134]^x[132]^x[130]^x[123]^x[118]^x[108]^x[106]^x[102]^x[97]^x[96]^x[89]^x[56]^x[46]^x[45]^x[44]^x[35]^x[34]^x[33]^x[8]^x[2];
	y[21]=x[375]^x[372]^x[365]^x[364]^x[362]^x[361]^x[354]^x[353]^x[346]^x[313]^x[311]^x[309]^x[307]^x[304]^x[302]^x[299]^x[296]^x[289]^x[288]^x[282]^x[277]^x[276]^x[271]^x[270]^x[267]^x[265]^x[259]^x[256]^x[242]^x[231]^x[220]^x[219]^x[218]^x[215]^x[213]^x[209]^x[208]^x[207]^x[205]^x[204]^x[203]^x[194]^x[193]^x[192]^x[182]^x[181]^x[171]^x[153]^x[151]^x[149]^x[145]^x[144]^x[143]^x[142]^x[138]^x[137]^x[132]^x[131]^x[129]^x[128]^x[122]^x[117]^x[107]^x[105]^x[101]^x[96]^x[88]^x[55]^x[45]^x[44]^x[43]^x[34]^x[33]^x[32]^x[7]^x[1];
	y[20]=x[383]^x[382]^x[374]^x[371]^x[364]^x[363]^x[360]^x[353]^x[352]^x[319]^x[318]^x[314]^x[313]^x[310]^x[308]^x[306]^x[302]^x[297]^x[288]^x[287]^x[281]^x[276]^x[275]^x[270]^x[269]^x[264]^x[258]^x[241]^x[230]^x[223]^x[219]^x[218]^x[217]^x[214]^x[212]^x[206]^x[204]^x[203]^x[197]^x[193]^x[192]^x[181]^x[180]^x[170]^x[159]^x[158]^x[154]^x[152]^x[150]^x[144]^x[142]^x[138]^x[137]^x[136]^x[132]^x[131]^x[130]^x[128]^x[127]^x[116]^x[115]^x[104]^x[66]^x[63]^x[54]^x[44]^x[43]^x[33]^x[32]^x[6]^x[0];
	y[19]=x[383]^x[382]^x[381]^x[373]^x[372]^x[371]^x[370]^x[363]^x[361]^x[359]^x[352]^x[319]^x[317]^x[309]^x[306]^x[305]^x[298]^x[296]^x[295]^x[286]^x[280]^x[275]^x[274]^x[269]^x[268]^x[263]^x[257]^x[240]^x[229]^x[223]^x[222]^x[218]^x[217]^x[216]^x[213]^x[211]^x[207]^x[205]^x[203]^x[192]^x[180]^x[179]^x[169]^x[159]^x[157]^x[153]^x[151]^x[149]^x[147]^x[143]^x[141]^x[138]^x[137]^x[136]^x[135]^x[132]^x[131]^x[130]^x[129]^x[126]^x[115]^x[114]^x[103]^x[63]^x[62]^x[53]^x[43]^x[32]^x[5];
	y[18]=x[383]^x[382]^x[381]^x[380]^x[372]^x[371]^x[370]^x[369]^x[360]^x[358]^x[318]^x[316]^x[308]^x[305]^x[304]^x[297]^x[295]^x[294]^x[285]^x[279]^x[274]^x[273]^x[268]^x[267]^x[262]^x[256]^x[239]^x[228]^x[223]^x[222]^x[221]^x[217]^x[216]^x[215]^x[212]^x[210]^x[206]^x[204]^x[179]^x[178]^x[168]^x[158]^x[156]^x[152]^x[150]^x[148]^x[146]^x[142]^x[140]^x[137]^x[136]^x[135]^x[134]^x[131]^x[130]^x[129]^x[128]^x[125]^x[114]^x[113]^x[102]^x[63]^x[62]^x[61]^x[52]^x[4];
	y[17]=x[382]^x[381]^x[380]^x[379]^x[371]^x[370]^x[369]^x[368]^x[359]^x[357]^x[317]^x[315]^x[310]^x[309]^x[307]^x[298]^x[296]^x[294]^x[292]^x[288]^x[284]^x[278]^x[273]^x[272]^x[267]^x[261]^x[238]^x[227]^x[222]^x[221]^x[220]^x[216]^x[215]^x[214]^x[211]^x[209]^x[205]^x[203]^x[178]^x[177]^x[167]^x[157]^x[155]^x[151]^x[150]^x[147]^x[145]^x[141]^x[139]^x[138]^x[136]^x[135]^x[134]^x[133]^x[130]^x[129]^x[124]^x[113]^x[112]^x[101]^x[62]^x[61]^x[60]^x[51]^x[3];
	y[16]=x[381]^x[380]^x[379]^x[378]^x[370]^x[369]^x[368]^x[367]^x[358]^x[356]^x[316]^x[314]^x[308]^x[306]^x[303]^x[297]^x[295]^x[293]^x[292]^x[291]^x[283]^x[277]^x[272]^x[271]^x[266]^x[260]^x[237]^x[226]^x[221]^x[220]^x[219]^x[215]^x[214]^x[213]^x[210]^x[208]^x[204]^x[202]^x[177]^x[176]^x[166]^x[156]^x[154]^x[150]^x[146]^x[144]^x[140]^x[138]^x[137]^x[135]^x[134]^x[133]^x[132]^x[129]^x[128]^x[123]^x[112]^x[111]^x[100]^x[61]^x[60]^x[59]^x[50]^x[2];
	y[15]=x[380]^x[379]^x[378]^x[377]^x[369]^x[368]^x[367]^x[366]^x[357]^x[355]^x[315]^x[313]^x[309]^x[307]^x[305]^x[303]^x[302]^x[298]^x[296]^x[294]^x[291]^x[290]^x[282]^x[276]^x[271]^x[270]^x[265]^x[259]^x[236]^x[225]^x[220]^x[219]^x[218]^x[214]^x[213]^x[212]^x[209]^x[207]^x[202]^x[201]^x[192]^x[176]^x[175]^x[165]^x[155]^x[153]^x[145]^x[143]^x[139]^x[138]^x[137]^x[136]^x[134]^x[133]^x[132]^x[131]^x[128]^x[122]^x[111]^x[110]^x[99]^x[60]^x[59]^x[58]^x[49]^x[1];
	y[14]=x[379]^x[378]^x[377]^x[376]^x[368]^x[367]^x[366]^x[365]^x[356]^x[354]^x[314]^x[312]^x[308]^x[306]^x[304]^x[302]^x[301]^x[297]^x[295]^x[293]^x[290]^x[289]^x[281]^x[275]^x[270]^x[269]^x[264]^x[258]^x[235]^x[224]^x[219]^x[218]^x[217]^x[213]^x[212]^x[211]^x[208]^x[206]^x[202]^x[201]^x[200]^x[175]^x[174]^x[164]^x[154]^x[152]^x[144]^x[142]^x[138]^x[137]^x[136]^x[135]^x[133]^x[132]^x[131]^x[130]^x[121]^x[110]^x[109]^x[98]^x[59]^x[58]^x[57]^x[48]^x[0];
	y[13]=x[378]^x[377]^x[376]^x[375]^x[367]^x[366]^x[365]^x[364]^x[355]^x[353]^x[313]^x[311]^x[307]^x[305]^x[303]^x[301]^x[300]^x[296]^x[294]^x[292]^x[289]^x[288]^x[280]^x[274]^x[269]^x[268]^x[263]^x[257]^x[218]^x[217]^x[216]^x[212]^x[211]^x[210]^x[207]^x[205]^x[201]^x[200]^x[199]^x[174]^x[173]^x[163]^x[153]^x[151]^x[143]^x[141]^x[137]^x[136]^x[135]^x[134]^x[132]^x[131]^x[130]^x[129]^x[120]^x[109]^x[108]^x[97]^x[58]^x[57]^x[56]^x[47];
	y[12]=x[377]^x[376]^x[375]^x[374]^x[366]^x[365]^x[364]^x[363]^x[354]^x[352]^x[312]^x[310]^x[306]^x[304]^x[302]^x[300]^x[295]^x[293]^x[291]^x[279]^x[273]^x[268]^x[267]^x[262]^x[256]^x[217]^x[216]^x[215]^x[211]^x[210]^x[209]^x[206]^x[204]^x[200]^x[199]^x[198]^x[173]^x[172]^x[162]^x[152]^x[150]^x[142]^x[140]^x[136]^x[135]^x[134]^x[133]^x[131]^x[130]^x[129]^x[128]^x[119]^x[108]^x[107]^x[96]^x[57]^x[56]^x[55]^x[46];
	y[11]=x[376]^x[375]^x[374]^x[365]^x[363]^x[352]^x[311]^x[310]^x[305]^x[304]^x[301]^x[294]^x[293]^x[290]^x[278]^x[272]^x[267]^x[261]^x[216]^x[215]^x[214]^x[210]^x[209]^x[208]^x[205]^x[203]^x[199]^x[198]^x[197]^x[172]^x[171]^x[161]^x[151]^x[150]^x[141]^x[135]^x[134]^x[133]^x[130]^x[129]^x[128]^x[118]^x[107]^x[56]^x[55]^x[54]^x[45];
	y[10]=x[375]^x[374]^x[373]^x[364]^x[363]^x[362]^x[352]^x[310]^x[304]^x[300]^x[298]^x[293]^x[289]^x[277]^x[271]^x[266]^x[260]^x[215]^x[214]^x[213]^x[209]^x[208]^x[207]^x[204]^x[202]^x[198]^x[197]^x[196]^x[171]^x[170]^x[160]^x[150]^x[140]^x[138]^x[134]^x[133]^x[132]^x[129]^x[128]^x[117]^x[106]^x[55]^x[54]^x[53]^x[44];
	y[9]=x[383]^x[382]^x[374]^x[373]^x[371]^x[363]^x[361]^x[317]^x[309]^x[308]^x[307]^x[299]^x[295]^x[288]^x[276]^x[270]^x[265]^x[259]^x[218]^x[214]^x[213]^x[212]^x[208]^x[207]^x[206]^x[203]^x[201]^x[197]^x[195]^x[191]^x[169]^x[149]^x[148]^x[147]^x[143]^x[142]^x[141]^x[139]^x[137]^x[133]^x[131]^x[128]^x[116]^x[105]^x[54]^x[53]^x[52]^x[43];
	y[8]=x[381]^x[373]^x[372]^x[371]^x[370]^x[362]^x[360]^x[319]^x[316]^x[308]^x[307]^x[306]^x[294]^x[275]^x[269]^x[264]^x[258]^x[213]^x[212]^x[211]^x[207]^x[206]^x[205]^x[202]^x[200]^x[196]^x[194]^x[190]^x[168]^x[159]^x[153]^x[148]^x[146]^x[142]^x[140]^x[136]^x[130]^x[115]^x[104]^x[53]^x[52]^x[51]^x[42];
	y[7]=x[380]^x[372]^x[371]^x[370]^x[369]^x[361]^x[359]^x[318]^x[315]^x[307]^x[306]^x[305]^x[293]^x[274]^x[268]^x[263]^x[257]^x[212]^x[211]^x[210]^x[206]^x[205]^x[204]^x[201]^x[199]^x[195]^x[193]^x[189]^x[167]^x[158]^x[152]^x[147]^x[145]^x[141]^x[139]^x[135]^x[129]^x[114]^x[103]^x[74]^x[52]^x[51]^x[50]^x[41];
	y[6]=x[379]^x[371]^x[370]^x[369]^x[368]^x[360]^x[358]^x[317]^x[314]^x[306]^x[305]^x[304]^x[292]^x[273]^x[267]^x[262]^x[256]^x[211]^x[210]^x[209]^x[205]^x[204]^x[203]^x[200]^x[198]^x[194]^x[192]^x[188]^x[166]^x[157]^x[151]^x[146]^x[144]^x[140]^x[138]^x[134]^x[128]^x[113]^x[102]^x[73]^x[51]^x[50]^x[49]^x[40];
	y[5]=x[378]^x[370]^x[369]^x[367]^x[359]^x[341]^x[330]^x[316]^x[313]^x[310]^x[305]^x[303]^x[293]^x[291]^x[288]^x[272]^x[261]^x[214]^x[210]^x[209]^x[208]^x[199]^x[197]^x[192]^x[187]^x[165]^x[156]^x[145]^x[143]^x[139]^x[137]^x[128]^x[112]^x[106]^x[101]^x[100]^x[72]^x[50]^x[49]^x[48]^x[39];
	y[4]=x[377]^x[369]^x[368]^x[367]^x[366]^x[358]^x[356]^x[340]^x[329]^x[315]^x[312]^x[309]^x[304]^x[302]^x[298]^x[292]^x[290]^x[271]^x[260]^x[209]^x[208]^x[207]^x[198]^x[196]^x[186]^x[164]^x[155]^x[144]^x[142]^x[136]^x[132]^x[111]^x[105]^x[100]^x[99]^x[71]^x[49]^x[48]^x[47]^x[38];
	y[3]=x[376]^x[368]^x[367]^x[366]^x[365]^x[357]^x[355]^x[339]^x[328]^x[314]^x[311]^x[308]^x[303]^x[301]^x[297]^x[291]^x[289]^x[270]^x[259]^x[208]^x[207]^x[206]^x[197]^x[195]^x[185]^x[163]^x[154]^x[143]^x[141]^x[135]^x[131]^x[110]^x[104]^x[99]^x[98]^x[70]^x[48]^x[47]^x[46]^x[37];
	y[2]=x[375]^x[367]^x[366]^x[365]^x[364]^x[356]^x[354]^x[338]^x[327]^x[313]^x[310]^x[307]^x[302]^x[300]^x[296]^x[290]^x[288]^x[269]^x[258]^x[207]^x[206]^x[205]^x[196]^x[194]^x[184]^x[162]^x[153]^x[142]^x[140]^x[134]^x[130]^x[109]^x[103]^x[98]^x[97]^x[69]^x[47]^x[46]^x[45]^x[36];
	y[1]=x[374]^x[366]^x[365]^x[364]^x[363]^x[355]^x[353]^x[337]^x[326]^x[312]^x[306]^x[301]^x[299]^x[295]^x[289]^x[268]^x[257]^x[206]^x[205]^x[204]^x[195]^x[193]^x[183]^x[161]^x[152]^x[141]^x[139]^x[133]^x[129]^x[108]^x[102]^x[97]^x[96]^x[46]^x[45]^x[44]^x[35];
	y[0]=x[374]^x[365]^x[364]^x[363]^x[354]^x[336]^x[325]^x[311]^x[305]^x[300]^x[299]^x[294]^x[267]^x[256]^x[205]^x[204]^x[203]^x[194]^x[192]^x[182]^x[160]^x[151]^x[140]^x[139]^x[133]^x[107]^x[101]^x[96]^x[45]^x[44]^x[43]^x[34];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint59(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[380]^x[374]^x[369]^x[363]^x[351]^x[350]^x[343]^x[342]^x[341]^x[340]^x[339]^x[331]^x[321]^x[282]^x[281]^x[277]^x[272]^x[270]^x[268]^x[267]^x[266]^x[263]^x[261]^x[257]^x[255]^x[254]^x[249]^x[248]^x[245]^x[243]^x[239]^x[237]^x[234]^x[228]^x[220]^x[209]^x[191]^x[187]^x[186]^x[185]^x[183]^x[182]^x[181]^x[177]^x[175]^x[171]^x[170]^x[166]^x[165]^x[164]^x[161]^x[159]^x[149]^x[145]^x[139]^x[133]^x[128]^x[122]^x[121]^x[117]^x[116]^x[115]^x[112]^x[111]^x[109]^x[108]^x[107]^x[102]^x[97]^x[96]^x[95]^x[94]^x[85]^x[83]^x[74]^x[34]^x[23]^x[22]^x[21]^x[11]^x[10]^x[7]^x[1];
	y[30]=x[379]^x[373]^x[368]^x[362]^x[350]^x[349]^x[342]^x[341]^x[340]^x[338]^x[330]^x[329]^x[320]^x[286]^x[285]^x[274]^x[267]^x[266]^x[262]^x[256]^x[254]^x[253]^x[248]^x[247]^x[244]^x[242]^x[238]^x[236]^x[233]^x[227]^x[219]^x[208]^x[190]^x[184]^x[182]^x[181]^x[180]^x[176]^x[175]^x[174]^x[170]^x[169]^x[165]^x[164]^x[163]^x[160]^x[159]^x[158]^x[148]^x[144]^x[132]^x[126]^x[120]^x[114]^x[108]^x[107]^x[106]^x[101]^x[100]^x[96]^x[94]^x[93]^x[84]^x[82]^x[73]^x[22]^x[21]^x[20]^x[10]^x[9]^x[6]^x[0];
	y[29]=x[378]^x[372]^x[367]^x[361]^x[351]^x[350]^x[349]^x[348]^x[341]^x[340]^x[337]^x[330]^x[329]^x[328]^x[287]^x[285]^x[284]^x[273]^x[265]^x[261]^x[253]^x[252]^x[247]^x[246]^x[243]^x[241]^x[237]^x[235]^x[232]^x[226]^x[218]^x[207]^x[191]^x[189]^x[185]^x[183]^x[181]^x[180]^x[179]^x[175]^x[174]^x[173]^x[170]^x[169]^x[168]^x[164]^x[163]^x[162]^x[158]^x[157]^x[147]^x[143]^x[131]^x[127]^x[125]^x[121]^x[119]^x[115]^x[113]^x[109]^x[107]^x[105]^x[99]^x[93]^x[92]^x[83]^x[81]^x[72]^x[43]^x[32]^x[31]^x[21]^x[20]^x[19]^x[10]^x[9]^x[8]^x[5];
	y[28]=x[377]^x[371]^x[366]^x[360]^x[350]^x[349]^x[348]^x[347]^x[340]^x[339]^x[336]^x[329]^x[328]^x[327]^x[286]^x[284]^x[283]^x[272]^x[264]^x[260]^x[252]^x[251]^x[246]^x[245]^x[242]^x[240]^x[236]^x[234]^x[231]^x[225]^x[217]^x[206]^x[190]^x[188]^x[184]^x[182]^x[180]^x[179]^x[178]^x[174]^x[173]^x[172]^x[169]^x[168]^x[167]^x[163]^x[162]^x[161]^x[157]^x[156]^x[146]^x[142]^x[130]^x[126]^x[124]^x[120]^x[118]^x[114]^x[112]^x[108]^x[106]^x[104]^x[98]^x[92]^x[91]^x[82]^x[80]^x[71]^x[42]^x[30]^x[20]^x[19]^x[18]^x[9]^x[8]^x[7]^x[4];
	y[27]=x[376]^x[370]^x[365]^x[359]^x[349]^x[348]^x[347]^x[346]^x[339]^x[338]^x[335]^x[328]^x[327]^x[326]^x[285]^x[283]^x[282]^x[271]^x[263]^x[259]^x[251]^x[250]^x[245]^x[244]^x[241]^x[239]^x[235]^x[233]^x[230]^x[224]^x[216]^x[205]^x[189]^x[187]^x[183]^x[181]^x[179]^x[178]^x[177]^x[173]^x[172]^x[171]^x[168]^x[167]^x[166]^x[162]^x[161]^x[160]^x[156]^x[155]^x[145]^x[141]^x[129]^x[125]^x[123]^x[119]^x[117]^x[113]^x[111]^x[107]^x[105]^x[103]^x[97]^x[91]^x[90]^x[81]^x[79]^x[70]^x[41]^x[29]^x[19]^x[18]^x[17]^x[8]^x[7]^x[6]^x[3];
	y[26]=x[375]^x[369]^x[364]^x[358]^x[348]^x[347]^x[345]^x[338]^x[337]^x[334]^x[327]^x[326]^x[325]^x[319]^x[287]^x[286]^x[284]^x[280]^x[277]^x[276]^x[275]^x[271]^x[269]^x[267]^x[262]^x[258]^x[256]^x[255]^x[250]^x[249]^x[244]^x[243]^x[240]^x[238]^x[232]^x[229]^x[215]^x[204]^x[191]^x[188]^x[186]^x[181]^x[180]^x[178]^x[177]^x[176]^x[172]^x[167]^x[166]^x[165]^x[161]^x[160]^x[155]^x[154]^x[144]^x[140]^x[128]^x[127]^x[126]^x[124]^x[118]^x[117]^x[116]^x[115]^x[112]^x[110]^x[107]^x[106]^x[104]^x[102]^x[101]^x[95]^x[90]^x[80]^x[78]^x[74]^x[69]^x[68]^x[61]^x[28]^x[18]^x[17]^x[16]^x[7]^x[6]^x[5]^x[2];
	y[25]=x[374]^x[368]^x[363]^x[357]^x[347]^x[346]^x[345]^x[344]^x[337]^x[336]^x[333]^x[326]^x[325]^x[324]^x[318]^x[285]^x[283]^x[281]^x[280]^x[279]^x[276]^x[274]^x[270]^x[269]^x[268]^x[261]^x[257]^x[254]^x[249]^x[248]^x[243]^x[242]^x[239]^x[237]^x[231]^x[228]^x[214]^x[203]^x[191]^x[190]^x[187]^x[185]^x[181]^x[180]^x[179]^x[177]^x[176]^x[175]^x[171]^x[166]^x[165]^x[164]^x[160]^x[154]^x[153]^x[143]^x[139]^x[125]^x[123]^x[121]^x[117]^x[116]^x[115]^x[114]^x[111]^x[109]^x[105]^x[103]^x[101]^x[94]^x[89]^x[79]^x[77]^x[73]^x[68]^x[67]^x[60]^x[39]^x[27]^x[17]^x[16]^x[15]^x[6]^x[5]^x[4]^x[1];
	y[24]=x[373]^x[367]^x[362]^x[356]^x[346]^x[345]^x[344]^x[343]^x[336]^x[335]^x[332]^x[325]^x[324]^x[323]^x[317]^x[284]^x[282]^x[280]^x[279]^x[278]^x[275]^x[273]^x[269]^x[268]^x[267]^x[260]^x[256]^x[253]^x[248]^x[247]^x[242]^x[241]^x[238]^x[236]^x[230]^x[227]^x[213]^x[202]^x[191]^x[190]^x[189]^x[186]^x[184]^x[180]^x[179]^x[178]^x[176]^x[175]^x[174]^x[165]^x[164]^x[163]^x[153]^x[152]^x[142]^x[138]^x[124]^x[122]^x[120]^x[116]^x[115]^x[114]^x[113]^x[110]^x[108]^x[104]^x[102]^x[100]^x[93]^x[88]^x[78]^x[76]^x[72]^x[67]^x[66]^x[59]^x[38]^x[26]^x[16]^x[15]^x[14]^x[5]^x[4]^x[3]^x[0];
	y[23]=x[372]^x[366]^x[361]^x[355]^x[345]^x[344]^x[343]^x[342]^x[335]^x[334]^x[331]^x[324]^x[323]^x[322]^x[316]^x[283]^x[281]^x[279]^x[277]^x[274]^x[272]^x[268]^x[266]^x[259]^x[252]^x[247]^x[246]^x[241]^x[240]^x[237]^x[235]^x[229]^x[226]^x[212]^x[201]^x[190]^x[189]^x[188]^x[185]^x[183]^x[179]^x[178]^x[177]^x[175]^x[174]^x[173]^x[164]^x[163]^x[162]^x[152]^x[151]^x[141]^x[137]^x[123]^x[121]^x[119]^x[115]^x[114]^x[113]^x[112]^x[109]^x[107]^x[103]^x[101]^x[99]^x[92]^x[87]^x[77]^x[75]^x[71]^x[66]^x[65]^x[58]^x[25]^x[15]^x[14]^x[13]^x[4]^x[3]^x[2];
	y[22]=x[371]^x[365]^x[360]^x[354]^x[344]^x[343]^x[342]^x[341]^x[334]^x[333]^x[330]^x[323]^x[322]^x[321]^x[315]^x[282]^x[280]^x[278]^x[276]^x[273]^x[271]^x[267]^x[265]^x[258]^x[251]^x[246]^x[245]^x[240]^x[239]^x[236]^x[234]^x[228]^x[225]^x[211]^x[200]^x[189]^x[188]^x[187]^x[184]^x[182]^x[178]^x[177]^x[176]^x[174]^x[173]^x[172]^x[163]^x[162]^x[161]^x[151]^x[150]^x[140]^x[136]^x[122]^x[120]^x[118]^x[114]^x[113]^x[112]^x[111]^x[108]^x[106]^x[102]^x[100]^x[98]^x[91]^x[86]^x[76]^x[74]^x[70]^x[65]^x[64]^x[57]^x[24]^x[14]^x[13]^x[12]^x[3]^x[2]^x[1];
	y[21]=x[370]^x[364]^x[359]^x[353]^x[343]^x[340]^x[333]^x[332]^x[330]^x[329]^x[322]^x[321]^x[314]^x[281]^x[279]^x[277]^x[275]^x[272]^x[270]^x[267]^x[264]^x[257]^x[256]^x[250]^x[245]^x[244]^x[239]^x[238]^x[235]^x[233]^x[227]^x[224]^x[210]^x[199]^x[188]^x[187]^x[186]^x[183]^x[181]^x[177]^x[176]^x[175]^x[173]^x[172]^x[171]^x[162]^x[161]^x[160]^x[150]^x[149]^x[139]^x[135]^x[121]^x[119]^x[117]^x[113]^x[112]^x[111]^x[110]^x[106]^x[105]^x[100]^x[99]^x[97]^x[96]^x[90]^x[85]^x[75]^x[73]^x[69]^x[64]^x[56]^x[23]^x[13]^x[12]^x[11]^x[2]^x[1]^x[0];
	y[20]=x[369]^x[363]^x[358]^x[352]^x[351]^x[350]^x[342]^x[339]^x[332]^x[331]^x[328]^x[321]^x[320]^x[287]^x[286]^x[282]^x[281]^x[278]^x[276]^x[274]^x[270]^x[265]^x[256]^x[255]^x[249]^x[244]^x[243]^x[238]^x[237]^x[232]^x[226]^x[209]^x[198]^x[191]^x[187]^x[186]^x[185]^x[182]^x[180]^x[174]^x[172]^x[171]^x[165]^x[161]^x[160]^x[149]^x[148]^x[138]^x[134]^x[127]^x[126]^x[122]^x[120]^x[118]^x[112]^x[110]^x[106]^x[105]^x[104]^x[100]^x[99]^x[98]^x[96]^x[95]^x[84]^x[83]^x[72]^x[34]^x[31]^x[22]^x[12]^x[11]^x[1]^x[0];
	y[19]=x[368]^x[357]^x[351]^x[350]^x[349]^x[341]^x[340]^x[339]^x[338]^x[331]^x[329]^x[327]^x[320]^x[287]^x[285]^x[277]^x[274]^x[273]^x[266]^x[264]^x[263]^x[254]^x[248]^x[243]^x[242]^x[237]^x[236]^x[231]^x[225]^x[208]^x[197]^x[191]^x[190]^x[186]^x[185]^x[184]^x[181]^x[179]^x[175]^x[173]^x[171]^x[160]^x[148]^x[147]^x[137]^x[133]^x[127]^x[125]^x[121]^x[119]^x[117]^x[115]^x[111]^x[109]^x[106]^x[105]^x[104]^x[103]^x[100]^x[99]^x[98]^x[97]^x[94]^x[83]^x[82]^x[71]^x[31]^x[30]^x[21]^x[11]^x[0];
	y[18]=x[367]^x[356]^x[351]^x[350]^x[349]^x[348]^x[340]^x[339]^x[338]^x[337]^x[328]^x[326]^x[286]^x[284]^x[276]^x[273]^x[272]^x[265]^x[263]^x[262]^x[253]^x[247]^x[242]^x[241]^x[236]^x[235]^x[230]^x[224]^x[207]^x[196]^x[191]^x[190]^x[189]^x[185]^x[184]^x[183]^x[180]^x[178]^x[174]^x[172]^x[147]^x[146]^x[136]^x[132]^x[126]^x[124]^x[120]^x[118]^x[116]^x[114]^x[110]^x[108]^x[105]^x[104]^x[103]^x[102]^x[99]^x[98]^x[97]^x[96]^x[93]^x[82]^x[81]^x[70]^x[31]^x[30]^x[29]^x[20];
	y[17]=x[366]^x[355]^x[350]^x[349]^x[348]^x[347]^x[339]^x[338]^x[337]^x[336]^x[327]^x[325]^x[285]^x[283]^x[278]^x[277]^x[275]^x[266]^x[264]^x[262]^x[260]^x[256]^x[252]^x[246]^x[241]^x[240]^x[235]^x[229]^x[206]^x[195]^x[190]^x[189]^x[188]^x[184]^x[183]^x[182]^x[179]^x[177]^x[173]^x[171]^x[146]^x[145]^x[135]^x[131]^x[125]^x[123]^x[119]^x[118]^x[115]^x[113]^x[109]^x[107]^x[106]^x[104]^x[103]^x[102]^x[101]^x[98]^x[97]^x[92]^x[81]^x[80]^x[69]^x[30]^x[29]^x[28]^x[19];
	y[16]=x[365]^x[354]^x[349]^x[348]^x[347]^x[346]^x[338]^x[337]^x[336]^x[335]^x[326]^x[324]^x[284]^x[282]^x[276]^x[274]^x[271]^x[265]^x[263]^x[261]^x[260]^x[259]^x[251]^x[245]^x[240]^x[239]^x[234]^x[228]^x[205]^x[194]^x[189]^x[188]^x[187]^x[183]^x[182]^x[181]^x[178]^x[176]^x[172]^x[170]^x[145]^x[144]^x[134]^x[130]^x[124]^x[122]^x[118]^x[114]^x[112]^x[108]^x[106]^x[105]^x[103]^x[102]^x[101]^x[100]^x[97]^x[96]^x[91]^x[80]^x[79]^x[68]^x[29]^x[28]^x[27]^x[18];
	y[15]=x[364]^x[353]^x[348]^x[347]^x[346]^x[345]^x[337]^x[336]^x[335]^x[334]^x[325]^x[323]^x[283]^x[281]^x[277]^x[275]^x[273]^x[271]^x[270]^x[266]^x[264]^x[262]^x[259]^x[258]^x[250]^x[244]^x[239]^x[238]^x[233]^x[227]^x[204]^x[193]^x[188]^x[187]^x[186]^x[182]^x[181]^x[180]^x[177]^x[175]^x[170]^x[169]^x[160]^x[144]^x[143]^x[133]^x[129]^x[123]^x[121]^x[113]^x[111]^x[107]^x[106]^x[105]^x[104]^x[102]^x[101]^x[100]^x[99]^x[96]^x[90]^x[79]^x[78]^x[67]^x[28]^x[27]^x[26]^x[17];
	y[14]=x[363]^x[352]^x[347]^x[346]^x[345]^x[344]^x[336]^x[335]^x[334]^x[333]^x[324]^x[322]^x[282]^x[280]^x[276]^x[274]^x[272]^x[270]^x[269]^x[265]^x[263]^x[261]^x[258]^x[257]^x[249]^x[243]^x[238]^x[237]^x[232]^x[226]^x[203]^x[192]^x[187]^x[186]^x[185]^x[181]^x[180]^x[179]^x[176]^x[174]^x[170]^x[169]^x[168]^x[143]^x[142]^x[132]^x[128]^x[122]^x[120]^x[112]^x[110]^x[106]^x[105]^x[104]^x[103]^x[101]^x[100]^x[99]^x[98]^x[89]^x[78]^x[77]^x[66]^x[27]^x[26]^x[25]^x[16];
	y[13]=x[346]^x[345]^x[344]^x[343]^x[335]^x[334]^x[333]^x[332]^x[323]^x[321]^x[281]^x[279]^x[275]^x[273]^x[271]^x[269]^x[268]^x[264]^x[262]^x[260]^x[257]^x[256]^x[248]^x[242]^x[237]^x[236]^x[231]^x[225]^x[186]^x[185]^x[184]^x[180]^x[179]^x[178]^x[175]^x[173]^x[169]^x[168]^x[167]^x[142]^x[141]^x[131]^x[121]^x[119]^x[111]^x[109]^x[105]^x[104]^x[103]^x[102]^x[100]^x[99]^x[98]^x[97]^x[88]^x[77]^x[76]^x[65]^x[26]^x[25]^x[24]^x[15];
	y[12]=x[345]^x[344]^x[343]^x[342]^x[334]^x[333]^x[332]^x[331]^x[322]^x[320]^x[280]^x[278]^x[274]^x[272]^x[270]^x[268]^x[263]^x[261]^x[259]^x[247]^x[241]^x[236]^x[235]^x[230]^x[224]^x[185]^x[184]^x[183]^x[179]^x[178]^x[177]^x[174]^x[172]^x[168]^x[167]^x[166]^x[141]^x[140]^x[130]^x[120]^x[118]^x[110]^x[108]^x[104]^x[103]^x[102]^x[101]^x[99]^x[98]^x[97]^x[96]^x[87]^x[76]^x[75]^x[64]^x[25]^x[24]^x[23]^x[14];
	y[11]=x[344]^x[343]^x[342]^x[333]^x[331]^x[320]^x[279]^x[278]^x[273]^x[272]^x[269]^x[262]^x[261]^x[258]^x[246]^x[240]^x[235]^x[229]^x[184]^x[183]^x[182]^x[178]^x[177]^x[176]^x[173]^x[171]^x[167]^x[166]^x[165]^x[140]^x[139]^x[129]^x[119]^x[118]^x[109]^x[103]^x[102]^x[101]^x[98]^x[97]^x[96]^x[86]^x[75]^x[24]^x[23]^x[22]^x[13];
	y[10]=x[343]^x[342]^x[341]^x[332]^x[331]^x[330]^x[320]^x[278]^x[272]^x[268]^x[266]^x[261]^x[257]^x[245]^x[239]^x[234]^x[228]^x[183]^x[182]^x[181]^x[177]^x[176]^x[175]^x[172]^x[170]^x[166]^x[165]^x[164]^x[139]^x[138]^x[128]^x[118]^x[108]^x[106]^x[102]^x[101]^x[100]^x[97]^x[96]^x[85]^x[74]^x[23]^x[22]^x[21]^x[12];
	y[9]=x[351]^x[350]^x[342]^x[341]^x[339]^x[331]^x[329]^x[285]^x[277]^x[276]^x[275]^x[267]^x[263]^x[256]^x[244]^x[238]^x[233]^x[227]^x[186]^x[182]^x[181]^x[180]^x[176]^x[175]^x[174]^x[171]^x[169]^x[165]^x[163]^x[159]^x[137]^x[117]^x[116]^x[115]^x[111]^x[110]^x[109]^x[107]^x[105]^x[101]^x[99]^x[96]^x[84]^x[73]^x[22]^x[21]^x[20]^x[11];
	y[8]=x[349]^x[341]^x[340]^x[339]^x[338]^x[330]^x[328]^x[287]^x[284]^x[276]^x[275]^x[274]^x[262]^x[243]^x[237]^x[232]^x[226]^x[181]^x[180]^x[179]^x[175]^x[174]^x[173]^x[170]^x[168]^x[164]^x[162]^x[158]^x[136]^x[127]^x[121]^x[116]^x[114]^x[110]^x[108]^x[104]^x[98]^x[83]^x[72]^x[21]^x[20]^x[19]^x[10];
	y[7]=x[348]^x[340]^x[339]^x[338]^x[337]^x[329]^x[327]^x[286]^x[283]^x[275]^x[274]^x[273]^x[261]^x[242]^x[236]^x[231]^x[225]^x[180]^x[179]^x[178]^x[174]^x[173]^x[172]^x[169]^x[167]^x[163]^x[161]^x[157]^x[135]^x[126]^x[120]^x[115]^x[113]^x[109]^x[107]^x[103]^x[97]^x[82]^x[71]^x[42]^x[20]^x[19]^x[18]^x[9];
	y[6]=x[347]^x[339]^x[338]^x[337]^x[336]^x[328]^x[326]^x[285]^x[282]^x[274]^x[273]^x[272]^x[260]^x[241]^x[235]^x[230]^x[224]^x[179]^x[178]^x[177]^x[173]^x[172]^x[171]^x[168]^x[166]^x[162]^x[160]^x[156]^x[134]^x[125]^x[119]^x[114]^x[112]^x[108]^x[106]^x[102]^x[96]^x[81]^x[70]^x[41]^x[19]^x[18]^x[17]^x[8];
	y[5]=x[346]^x[338]^x[337]^x[335]^x[327]^x[309]^x[298]^x[284]^x[281]^x[278]^x[273]^x[271]^x[261]^x[259]^x[256]^x[240]^x[229]^x[182]^x[178]^x[177]^x[176]^x[167]^x[165]^x[160]^x[155]^x[133]^x[124]^x[113]^x[111]^x[107]^x[105]^x[96]^x[80]^x[74]^x[69]^x[68]^x[40]^x[18]^x[17]^x[16]^x[7];
	y[4]=x[345]^x[337]^x[336]^x[335]^x[334]^x[326]^x[324]^x[308]^x[297]^x[283]^x[280]^x[277]^x[272]^x[270]^x[266]^x[260]^x[258]^x[239]^x[228]^x[177]^x[176]^x[175]^x[166]^x[164]^x[154]^x[132]^x[123]^x[112]^x[110]^x[104]^x[100]^x[79]^x[73]^x[68]^x[67]^x[39]^x[17]^x[16]^x[15]^x[6];
	y[3]=x[344]^x[336]^x[335]^x[334]^x[333]^x[325]^x[323]^x[307]^x[296]^x[282]^x[279]^x[276]^x[271]^x[269]^x[265]^x[259]^x[257]^x[238]^x[227]^x[176]^x[175]^x[174]^x[165]^x[163]^x[153]^x[131]^x[122]^x[111]^x[109]^x[103]^x[99]^x[78]^x[72]^x[67]^x[66]^x[38]^x[16]^x[15]^x[14]^x[5];
	y[2]=x[343]^x[335]^x[334]^x[333]^x[332]^x[324]^x[322]^x[306]^x[295]^x[281]^x[278]^x[275]^x[270]^x[268]^x[264]^x[258]^x[256]^x[237]^x[226]^x[175]^x[174]^x[173]^x[164]^x[162]^x[152]^x[130]^x[121]^x[110]^x[108]^x[102]^x[98]^x[77]^x[71]^x[66]^x[65]^x[37]^x[15]^x[14]^x[13]^x[4];
	y[1]=x[342]^x[334]^x[333]^x[332]^x[331]^x[323]^x[321]^x[305]^x[294]^x[280]^x[274]^x[269]^x[267]^x[263]^x[257]^x[236]^x[225]^x[174]^x[173]^x[172]^x[163]^x[161]^x[151]^x[129]^x[120]^x[109]^x[107]^x[101]^x[97]^x[76]^x[70]^x[65]^x[64]^x[14]^x[13]^x[12]^x[3];
	y[0]=x[342]^x[333]^x[332]^x[331]^x[322]^x[304]^x[293]^x[279]^x[273]^x[268]^x[267]^x[262]^x[235]^x[224]^x[173]^x[172]^x[171]^x[162]^x[160]^x[150]^x[128]^x[119]^x[108]^x[107]^x[101]^x[75]^x[69]^x[64]^x[13]^x[12]^x[11]^x[2];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint60(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[375]^x[370]^x[365]^x[362]^x[359]^x[354]^x[352]^x[348]^x[342]^x[337]^x[331]^x[319]^x[318]^x[311]^x[310]^x[309]^x[308]^x[307]^x[299]^x[289]^x[250]^x[249]^x[245]^x[240]^x[238]^x[236]^x[235]^x[234]^x[231]^x[229]^x[225]^x[223]^x[222]^x[217]^x[216]^x[213]^x[211]^x[207]^x[205]^x[202]^x[196]^x[188]^x[177]^x[159]^x[155]^x[154]^x[153]^x[144]^x[135]^x[134]^x[129]^x[127]^x[117]^x[113]^x[107]^x[101]^x[96]^x[90]^x[89]^x[85]^x[84]^x[83]^x[80]^x[79]^x[77]^x[76]^x[75]^x[70]^x[65]^x[64]^x[63]^x[62]^x[53]^x[51]^x[42]^x[2];
	y[30]=x[383]^x[374]^x[369]^x[364]^x[362]^x[361]^x[358]^x[353]^x[347]^x[341]^x[336]^x[330]^x[318]^x[317]^x[310]^x[309]^x[308]^x[306]^x[298]^x[297]^x[288]^x[254]^x[253]^x[242]^x[235]^x[234]^x[230]^x[224]^x[222]^x[221]^x[216]^x[215]^x[212]^x[210]^x[206]^x[204]^x[201]^x[195]^x[187]^x[176]^x[158]^x[152]^x[134]^x[133]^x[128]^x[127]^x[126]^x[116]^x[112]^x[100]^x[94]^x[88]^x[82]^x[76]^x[75]^x[74]^x[69]^x[68]^x[64]^x[62]^x[61]^x[52]^x[50]^x[41];
	y[29]=x[382]^x[373]^x[368]^x[363]^x[361]^x[360]^x[357]^x[352]^x[346]^x[340]^x[335]^x[329]^x[319]^x[318]^x[317]^x[316]^x[309]^x[308]^x[305]^x[298]^x[297]^x[296]^x[255]^x[253]^x[252]^x[241]^x[233]^x[229]^x[221]^x[220]^x[215]^x[214]^x[211]^x[209]^x[205]^x[203]^x[200]^x[194]^x[186]^x[175]^x[157]^x[151]^x[133]^x[126]^x[125]^x[115]^x[111]^x[99]^x[95]^x[93]^x[89]^x[87]^x[83]^x[81]^x[77]^x[75]^x[73]^x[67]^x[61]^x[60]^x[51]^x[49]^x[40]^x[11]^x[0];
	y[28]=x[383]^x[381]^x[372]^x[367]^x[360]^x[359]^x[356]^x[345]^x[339]^x[334]^x[328]^x[318]^x[317]^x[316]^x[315]^x[308]^x[307]^x[304]^x[297]^x[296]^x[295]^x[254]^x[252]^x[251]^x[240]^x[232]^x[228]^x[220]^x[219]^x[214]^x[213]^x[210]^x[208]^x[204]^x[202]^x[199]^x[193]^x[185]^x[174]^x[156]^x[150]^x[132]^x[125]^x[124]^x[114]^x[110]^x[98]^x[94]^x[92]^x[88]^x[86]^x[82]^x[80]^x[76]^x[74]^x[72]^x[66]^x[60]^x[59]^x[50]^x[48]^x[39]^x[10];
	y[27]=x[382]^x[380]^x[371]^x[366]^x[359]^x[358]^x[355]^x[344]^x[338]^x[333]^x[327]^x[317]^x[316]^x[315]^x[314]^x[307]^x[306]^x[303]^x[296]^x[295]^x[294]^x[253]^x[251]^x[250]^x[239]^x[231]^x[227]^x[219]^x[218]^x[213]^x[212]^x[209]^x[207]^x[203]^x[201]^x[198]^x[192]^x[184]^x[173]^x[155]^x[149]^x[131]^x[124]^x[123]^x[113]^x[109]^x[97]^x[93]^x[91]^x[87]^x[85]^x[81]^x[79]^x[75]^x[73]^x[71]^x[65]^x[59]^x[58]^x[49]^x[47]^x[38]^x[9];
	y[26]=x[381]^x[379]^x[370]^x[365]^x[358]^x[357]^x[354]^x[343]^x[337]^x[332]^x[326]^x[316]^x[315]^x[313]^x[306]^x[305]^x[302]^x[295]^x[294]^x[293]^x[287]^x[255]^x[254]^x[252]^x[248]^x[245]^x[244]^x[243]^x[239]^x[237]^x[235]^x[230]^x[226]^x[224]^x[223]^x[218]^x[217]^x[212]^x[211]^x[208]^x[206]^x[200]^x[197]^x[183]^x[172]^x[159]^x[154]^x[150]^x[149]^x[148]^x[139]^x[138]^x[130]^x[123]^x[122]^x[112]^x[108]^x[96]^x[95]^x[94]^x[92]^x[86]^x[85]^x[84]^x[83]^x[80]^x[78]^x[75]^x[74]^x[72]^x[70]^x[69]^x[63]^x[58]^x[48]^x[46]^x[42]^x[37]^x[36]^x[29];
	y[25]=x[380]^x[378]^x[369]^x[364]^x[357]^x[356]^x[353]^x[342]^x[336]^x[331]^x[325]^x[315]^x[314]^x[313]^x[312]^x[305]^x[304]^x[301]^x[294]^x[293]^x[292]^x[286]^x[253]^x[251]^x[249]^x[248]^x[247]^x[244]^x[242]^x[238]^x[237]^x[236]^x[229]^x[225]^x[222]^x[217]^x[216]^x[211]^x[210]^x[207]^x[205]^x[199]^x[196]^x[182]^x[171]^x[159]^x[158]^x[153]^x[148]^x[147]^x[138]^x[137]^x[129]^x[122]^x[121]^x[111]^x[107]^x[93]^x[91]^x[89]^x[85]^x[84]^x[83]^x[82]^x[79]^x[77]^x[73]^x[71]^x[69]^x[62]^x[57]^x[47]^x[45]^x[41]^x[36]^x[35]^x[28]^x[7];
	y[24]=x[379]^x[377]^x[368]^x[363]^x[356]^x[355]^x[352]^x[341]^x[335]^x[330]^x[324]^x[314]^x[313]^x[312]^x[311]^x[304]^x[303]^x[300]^x[293]^x[292]^x[291]^x[285]^x[252]^x[250]^x[248]^x[247]^x[246]^x[243]^x[241]^x[237]^x[236]^x[235]^x[228]^x[224]^x[221]^x[216]^x[215]^x[210]^x[209]^x[206]^x[204]^x[198]^x[195]^x[181]^x[170]^x[159]^x[158]^x[157]^x[152]^x[147]^x[146]^x[138]^x[137]^x[136]^x[128]^x[121]^x[120]^x[110]^x[106]^x[92]^x[90]^x[88]^x[84]^x[83]^x[82]^x[81]^x[78]^x[76]^x[72]^x[70]^x[68]^x[61]^x[56]^x[46]^x[44]^x[40]^x[35]^x[34]^x[27]^x[6];
	y[23]=x[378]^x[376]^x[367]^x[355]^x[354]^x[340]^x[334]^x[329]^x[323]^x[313]^x[312]^x[311]^x[310]^x[303]^x[302]^x[299]^x[292]^x[291]^x[290]^x[284]^x[251]^x[249]^x[247]^x[245]^x[242]^x[240]^x[236]^x[234]^x[227]^x[220]^x[215]^x[214]^x[209]^x[208]^x[205]^x[203]^x[197]^x[194]^x[180]^x[169]^x[158]^x[157]^x[156]^x[151]^x[146]^x[145]^x[137]^x[136]^x[135]^x[120]^x[119]^x[109]^x[105]^x[91]^x[89]^x[87]^x[83]^x[82]^x[81]^x[80]^x[77]^x[75]^x[71]^x[69]^x[67]^x[60]^x[55]^x[45]^x[43]^x[39]^x[34]^x[33]^x[26];
	y[22]=x[377]^x[375]^x[366]^x[354]^x[353]^x[339]^x[333]^x[328]^x[322]^x[312]^x[311]^x[310]^x[309]^x[302]^x[301]^x[298]^x[291]^x[290]^x[289]^x[283]^x[250]^x[248]^x[246]^x[244]^x[241]^x[239]^x[235]^x[233]^x[226]^x[219]^x[214]^x[213]^x[208]^x[207]^x[204]^x[202]^x[196]^x[193]^x[179]^x[168]^x[157]^x[156]^x[155]^x[150]^x[145]^x[144]^x[136]^x[135]^x[134]^x[119]^x[118]^x[108]^x[104]^x[90]^x[88]^x[86]^x[82]^x[81]^x[80]^x[79]^x[76]^x[74]^x[70]^x[68]^x[66]^x[59]^x[54]^x[44]^x[42]^x[38]^x[33]^x[32]^x[25];
	y[21]=x[376]^x[374]^x[365]^x[353]^x[352]^x[338]^x[332]^x[327]^x[321]^x[311]^x[308]^x[301]^x[300]^x[298]^x[297]^x[290]^x[289]^x[282]^x[249]^x[247]^x[245]^x[243]^x[240]^x[238]^x[235]^x[232]^x[225]^x[224]^x[218]^x[213]^x[212]^x[207]^x[206]^x[203]^x[201]^x[195]^x[192]^x[178]^x[167]^x[156]^x[155]^x[154]^x[149]^x[144]^x[143]^x[135]^x[134]^x[133]^x[118]^x[117]^x[107]^x[103]^x[89]^x[87]^x[85]^x[81]^x[80]^x[79]^x[78]^x[74]^x[73]^x[68]^x[67]^x[65]^x[64]^x[58]^x[53]^x[43]^x[41]^x[37]^x[32]^x[24];
	y[20]=x[383]^x[375]^x[373]^x[364]^x[362]^x[352]^x[337]^x[331]^x[326]^x[320]^x[319]^x[318]^x[310]^x[307]^x[300]^x[299]^x[296]^x[289]^x[288]^x[255]^x[254]^x[250]^x[249]^x[246]^x[244]^x[242]^x[238]^x[233]^x[224]^x[223]^x[217]^x[212]^x[211]^x[206]^x[205]^x[200]^x[194]^x[177]^x[166]^x[155]^x[154]^x[148]^x[144]^x[142]^x[134]^x[117]^x[116]^x[106]^x[102]^x[95]^x[94]^x[90]^x[88]^x[86]^x[80]^x[78]^x[74]^x[73]^x[72]^x[68]^x[67]^x[66]^x[64]^x[63]^x[52]^x[51]^x[40]^x[2];
	y[19]=x[383]^x[382]^x[374]^x[372]^x[363]^x[362]^x[361]^x[336]^x[325]^x[319]^x[318]^x[317]^x[309]^x[308]^x[307]^x[306]^x[299]^x[297]^x[295]^x[288]^x[255]^x[253]^x[245]^x[242]^x[241]^x[234]^x[232]^x[231]^x[222]^x[216]^x[211]^x[210]^x[205]^x[204]^x[199]^x[193]^x[176]^x[165]^x[154]^x[147]^x[141]^x[133]^x[116]^x[115]^x[105]^x[101]^x[95]^x[93]^x[89]^x[87]^x[85]^x[83]^x[79]^x[77]^x[74]^x[73]^x[72]^x[71]^x[68]^x[67]^x[66]^x[65]^x[62]^x[51]^x[50]^x[39];
	y[18]=x[382]^x[381]^x[373]^x[371]^x[362]^x[361]^x[360]^x[335]^x[324]^x[319]^x[318]^x[317]^x[316]^x[308]^x[307]^x[306]^x[305]^x[296]^x[294]^x[254]^x[252]^x[244]^x[241]^x[240]^x[233]^x[231]^x[230]^x[221]^x[215]^x[210]^x[209]^x[204]^x[203]^x[198]^x[192]^x[175]^x[164]^x[146]^x[140]^x[115]^x[114]^x[104]^x[100]^x[94]^x[92]^x[88]^x[86]^x[84]^x[82]^x[78]^x[76]^x[73]^x[72]^x[71]^x[70]^x[67]^x[66]^x[65]^x[64]^x[61]^x[50]^x[49]^x[38];
	y[17]=x[381]^x[380]^x[372]^x[370]^x[361]^x[360]^x[359]^x[334]^x[323]^x[318]^x[317]^x[316]^x[315]^x[307]^x[306]^x[305]^x[304]^x[295]^x[293]^x[253]^x[251]^x[246]^x[245]^x[243]^x[234]^x[232]^x[230]^x[228]^x[224]^x[220]^x[214]^x[209]^x[208]^x[203]^x[197]^x[174]^x[163]^x[145]^x[139]^x[114]^x[113]^x[103]^x[99]^x[93]^x[91]^x[87]^x[86]^x[83]^x[81]^x[77]^x[75]^x[74]^x[72]^x[71]^x[70]^x[69]^x[66]^x[65]^x[60]^x[49]^x[48]^x[37];
	y[16]=x[380]^x[379]^x[371]^x[369]^x[360]^x[359]^x[358]^x[333]^x[322]^x[317]^x[316]^x[315]^x[314]^x[306]^x[305]^x[304]^x[303]^x[294]^x[292]^x[252]^x[250]^x[244]^x[242]^x[239]^x[233]^x[231]^x[229]^x[228]^x[227]^x[219]^x[213]^x[208]^x[207]^x[202]^x[196]^x[173]^x[162]^x[144]^x[138]^x[113]^x[112]^x[102]^x[98]^x[92]^x[90]^x[86]^x[82]^x[80]^x[76]^x[74]^x[73]^x[71]^x[70]^x[69]^x[68]^x[65]^x[64]^x[59]^x[48]^x[47]^x[36];
	y[15]=x[379]^x[378]^x[370]^x[368]^x[359]^x[358]^x[357]^x[332]^x[321]^x[316]^x[315]^x[314]^x[313]^x[305]^x[304]^x[303]^x[302]^x[293]^x[291]^x[251]^x[249]^x[245]^x[243]^x[241]^x[239]^x[238]^x[234]^x[232]^x[230]^x[227]^x[226]^x[218]^x[212]^x[207]^x[206]^x[201]^x[195]^x[172]^x[161]^x[143]^x[139]^x[138]^x[137]^x[128]^x[112]^x[111]^x[101]^x[97]^x[91]^x[89]^x[81]^x[79]^x[75]^x[74]^x[73]^x[72]^x[70]^x[69]^x[68]^x[67]^x[64]^x[58]^x[47]^x[46]^x[35];
	y[14]=x[378]^x[377]^x[369]^x[367]^x[358]^x[357]^x[356]^x[331]^x[320]^x[315]^x[314]^x[313]^x[312]^x[304]^x[303]^x[302]^x[301]^x[292]^x[290]^x[250]^x[248]^x[244]^x[242]^x[240]^x[238]^x[237]^x[233]^x[231]^x[229]^x[226]^x[225]^x[217]^x[211]^x[206]^x[205]^x[200]^x[194]^x[171]^x[160]^x[142]^x[137]^x[136]^x[111]^x[110]^x[100]^x[96]^x[90]^x[88]^x[80]^x[78]^x[74]^x[73]^x[72]^x[71]^x[69]^x[68]^x[67]^x[66]^x[57]^x[46]^x[45]^x[34];
	y[13]=x[377]^x[376]^x[368]^x[366]^x[357]^x[356]^x[355]^x[314]^x[313]^x[312]^x[311]^x[303]^x[302]^x[301]^x[300]^x[291]^x[289]^x[249]^x[247]^x[243]^x[241]^x[239]^x[237]^x[236]^x[232]^x[230]^x[228]^x[225]^x[224]^x[216]^x[210]^x[205]^x[204]^x[199]^x[193]^x[141]^x[136]^x[135]^x[110]^x[109]^x[99]^x[89]^x[87]^x[79]^x[77]^x[73]^x[72]^x[71]^x[70]^x[68]^x[67]^x[66]^x[65]^x[56]^x[45]^x[44]^x[33];
	y[12]=x[376]^x[375]^x[367]^x[365]^x[356]^x[355]^x[354]^x[313]^x[312]^x[311]^x[310]^x[302]^x[301]^x[300]^x[299]^x[290]^x[288]^x[248]^x[246]^x[242]^x[240]^x[238]^x[236]^x[231]^x[229]^x[227]^x[215]^x[209]^x[204]^x[203]^x[198]^x[192]^x[140]^x[135]^x[134]^x[109]^x[108]^x[98]^x[88]^x[86]^x[78]^x[76]^x[72]^x[71]^x[70]^x[69]^x[67]^x[66]^x[65]^x[64]^x[55]^x[44]^x[43]^x[32];
	y[11]=x[375]^x[374]^x[366]^x[364]^x[355]^x[354]^x[353]^x[312]^x[311]^x[310]^x[301]^x[299]^x[288]^x[247]^x[246]^x[241]^x[240]^x[237]^x[230]^x[229]^x[226]^x[214]^x[208]^x[203]^x[197]^x[139]^x[134]^x[133]^x[108]^x[107]^x[97]^x[87]^x[86]^x[77]^x[71]^x[70]^x[69]^x[66]^x[65]^x[64]^x[54]^x[43];
	y[10]=x[374]^x[373]^x[365]^x[363]^x[354]^x[353]^x[352]^x[311]^x[310]^x[309]^x[300]^x[299]^x[298]^x[288]^x[246]^x[240]^x[236]^x[234]^x[229]^x[225]^x[213]^x[207]^x[202]^x[196]^x[138]^x[133]^x[132]^x[107]^x[106]^x[96]^x[86]^x[76]^x[74]^x[70]^x[69]^x[68]^x[65]^x[64]^x[53]^x[42];
	y[9]=x[383]^x[373]^x[372]^x[364]^x[353]^x[352]^x[319]^x[318]^x[310]^x[309]^x[307]^x[299]^x[297]^x[253]^x[245]^x[244]^x[243]^x[235]^x[231]^x[224]^x[212]^x[206]^x[201]^x[195]^x[154]^x[137]^x[131]^x[127]^x[105]^x[85]^x[84]^x[83]^x[79]^x[78]^x[77]^x[75]^x[73]^x[69]^x[67]^x[64]^x[52]^x[41];
	y[8]=x[383]^x[382]^x[372]^x[371]^x[363]^x[362]^x[352]^x[317]^x[309]^x[308]^x[307]^x[306]^x[298]^x[296]^x[255]^x[252]^x[244]^x[243]^x[242]^x[230]^x[211]^x[205]^x[200]^x[194]^x[136]^x[130]^x[126]^x[104]^x[95]^x[89]^x[84]^x[82]^x[78]^x[76]^x[72]^x[66]^x[51]^x[40];
	y[7]=x[383]^x[382]^x[381]^x[371]^x[370]^x[361]^x[316]^x[308]^x[307]^x[306]^x[305]^x[297]^x[295]^x[254]^x[251]^x[243]^x[242]^x[241]^x[229]^x[210]^x[204]^x[199]^x[193]^x[135]^x[129]^x[125]^x[103]^x[94]^x[88]^x[83]^x[81]^x[77]^x[75]^x[71]^x[65]^x[50]^x[39]^x[10];
	y[6]=x[382]^x[381]^x[380]^x[370]^x[369]^x[360]^x[315]^x[307]^x[306]^x[305]^x[304]^x[296]^x[294]^x[253]^x[250]^x[242]^x[241]^x[240]^x[228]^x[209]^x[203]^x[198]^x[192]^x[134]^x[128]^x[124]^x[102]^x[93]^x[87]^x[82]^x[80]^x[76]^x[74]^x[70]^x[64]^x[49]^x[38]^x[9];
	y[5]=x[381]^x[380]^x[379]^x[369]^x[368]^x[359]^x[314]^x[306]^x[305]^x[303]^x[295]^x[277]^x[266]^x[252]^x[249]^x[246]^x[241]^x[239]^x[229]^x[227]^x[224]^x[208]^x[197]^x[150]^x[140]^x[139]^x[138]^x[133]^x[129]^x[128]^x[123]^x[101]^x[92]^x[81]^x[79]^x[75]^x[73]^x[64]^x[48]^x[42]^x[37]^x[36]^x[8];
	y[4]=x[380]^x[379]^x[378]^x[368]^x[367]^x[358]^x[313]^x[305]^x[304]^x[303]^x[302]^x[294]^x[292]^x[276]^x[265]^x[251]^x[248]^x[245]^x[240]^x[238]^x[234]^x[228]^x[226]^x[207]^x[196]^x[139]^x[138]^x[137]^x[132]^x[128]^x[122]^x[100]^x[91]^x[80]^x[78]^x[72]^x[68]^x[47]^x[41]^x[36]^x[35]^x[7];
	y[3]=x[379]^x[378]^x[377]^x[367]^x[366]^x[357]^x[312]^x[304]^x[303]^x[302]^x[301]^x[293]^x[291]^x[275]^x[264]^x[250]^x[247]^x[244]^x[239]^x[237]^x[233]^x[227]^x[225]^x[206]^x[195]^x[138]^x[137]^x[136]^x[131]^x[121]^x[99]^x[90]^x[79]^x[77]^x[71]^x[67]^x[46]^x[40]^x[35]^x[34]^x[6];
	y[2]=x[378]^x[377]^x[376]^x[366]^x[365]^x[356]^x[311]^x[303]^x[302]^x[301]^x[300]^x[292]^x[290]^x[274]^x[263]^x[249]^x[246]^x[243]^x[238]^x[236]^x[232]^x[226]^x[224]^x[205]^x[194]^x[137]^x[136]^x[135]^x[130]^x[120]^x[98]^x[89]^x[78]^x[76]^x[70]^x[66]^x[45]^x[39]^x[34]^x[33]^x[5];
	y[1]=x[377]^x[376]^x[375]^x[365]^x[364]^x[355]^x[310]^x[302]^x[301]^x[300]^x[299]^x[291]^x[289]^x[273]^x[262]^x[248]^x[242]^x[237]^x[235]^x[231]^x[225]^x[204]^x[193]^x[136]^x[135]^x[134]^x[129]^x[119]^x[97]^x[88]^x[77]^x[75]^x[69]^x[65]^x[44]^x[38]^x[33]^x[32];
	y[0]=x[376]^x[375]^x[374]^x[364]^x[363]^x[354]^x[310]^x[301]^x[300]^x[299]^x[290]^x[272]^x[261]^x[247]^x[241]^x[236]^x[235]^x[230]^x[203]^x[192]^x[135]^x[134]^x[133]^x[128]^x[118]^x[96]^x[87]^x[76]^x[75]^x[69]^x[43]^x[37]^x[32];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint61(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[365]^x[354]^x[343]^x[338]^x[333]^x[330]^x[327]^x[322]^x[320]^x[316]^x[310]^x[305]^x[299]^x[287]^x[286]^x[279]^x[278]^x[277]^x[276]^x[275]^x[267]^x[257]^x[218]^x[217]^x[213]^x[208]^x[206]^x[204]^x[203]^x[202]^x[199]^x[197]^x[193]^x[191]^x[190]^x[185]^x[184]^x[181]^x[179]^x[175]^x[173]^x[170]^x[164]^x[156]^x[145]^x[130]^x[127]^x[123]^x[122]^x[121]^x[112]^x[103]^x[102]^x[97]^x[95]^x[85]^x[81]^x[75]^x[69]^x[64]^x[58]^x[57]^x[53]^x[52]^x[51]^x[48]^x[47]^x[45]^x[44]^x[43]^x[38]^x[33]^x[32]^x[31]^x[30]^x[21]^x[19]^x[10];
	y[30]=x[351]^x[342]^x[337]^x[332]^x[330]^x[329]^x[326]^x[321]^x[315]^x[309]^x[304]^x[298]^x[286]^x[285]^x[278]^x[277]^x[276]^x[274]^x[266]^x[265]^x[256]^x[222]^x[221]^x[210]^x[203]^x[202]^x[198]^x[192]^x[190]^x[189]^x[184]^x[183]^x[180]^x[178]^x[174]^x[172]^x[169]^x[163]^x[155]^x[144]^x[126]^x[120]^x[102]^x[101]^x[96]^x[95]^x[94]^x[84]^x[80]^x[68]^x[62]^x[56]^x[50]^x[44]^x[43]^x[42]^x[37]^x[36]^x[32]^x[30]^x[29]^x[20]^x[18]^x[9];
	y[29]=x[374]^x[352]^x[350]^x[341]^x[336]^x[331]^x[329]^x[328]^x[325]^x[320]^x[314]^x[308]^x[303]^x[297]^x[287]^x[286]^x[285]^x[284]^x[277]^x[276]^x[273]^x[266]^x[265]^x[264]^x[223]^x[221]^x[220]^x[209]^x[201]^x[197]^x[189]^x[188]^x[183]^x[182]^x[179]^x[177]^x[173]^x[171]^x[168]^x[162]^x[154]^x[143]^x[139]^x[133]^x[128]^x[125]^x[119]^x[101]^x[94]^x[93]^x[83]^x[79]^x[67]^x[63]^x[61]^x[57]^x[55]^x[51]^x[49]^x[45]^x[43]^x[41]^x[35]^x[29]^x[28]^x[19]^x[17]^x[8];
	y[28]=x[373]^x[362]^x[351]^x[349]^x[340]^x[335]^x[328]^x[327]^x[324]^x[313]^x[307]^x[302]^x[296]^x[286]^x[285]^x[284]^x[283]^x[276]^x[275]^x[272]^x[265]^x[264]^x[263]^x[222]^x[220]^x[219]^x[208]^x[200]^x[196]^x[188]^x[187]^x[182]^x[181]^x[178]^x[176]^x[172]^x[170]^x[167]^x[161]^x[153]^x[142]^x[138]^x[132]^x[124]^x[118]^x[100]^x[93]^x[92]^x[82]^x[78]^x[66]^x[62]^x[60]^x[56]^x[54]^x[50]^x[48]^x[44]^x[42]^x[40]^x[34]^x[28]^x[27]^x[18]^x[16]^x[7];
	y[27]=x[372]^x[361]^x[350]^x[348]^x[339]^x[334]^x[327]^x[326]^x[323]^x[312]^x[306]^x[301]^x[295]^x[285]^x[284]^x[283]^x[282]^x[275]^x[274]^x[271]^x[264]^x[263]^x[262]^x[221]^x[219]^x[218]^x[207]^x[199]^x[195]^x[187]^x[186]^x[181]^x[180]^x[177]^x[175]^x[171]^x[169]^x[166]^x[160]^x[152]^x[141]^x[137]^x[131]^x[123]^x[117]^x[99]^x[92]^x[91]^x[81]^x[77]^x[65]^x[61]^x[59]^x[55]^x[53]^x[49]^x[47]^x[43]^x[41]^x[39]^x[33]^x[27]^x[26]^x[17]^x[15]^x[6];
	y[26]=x[381]^x[371]^x[360]^x[349]^x[347]^x[338]^x[333]^x[326]^x[325]^x[322]^x[311]^x[305]^x[300]^x[294]^x[284]^x[283]^x[281]^x[274]^x[273]^x[270]^x[263]^x[262]^x[261]^x[255]^x[223]^x[222]^x[220]^x[216]^x[213]^x[212]^x[211]^x[207]^x[205]^x[203]^x[198]^x[194]^x[192]^x[191]^x[186]^x[185]^x[180]^x[179]^x[176]^x[174]^x[168]^x[165]^x[157]^x[140]^x[127]^x[122]^x[118]^x[117]^x[116]^x[107]^x[106]^x[98]^x[91]^x[90]^x[80]^x[76]^x[64]^x[63]^x[62]^x[60]^x[54]^x[53]^x[52]^x[51]^x[48]^x[46]^x[43]^x[42]^x[40]^x[38]^x[37]^x[31]^x[26]^x[16]^x[14]^x[10]^x[5]^x[4];
	y[25]=x[380]^x[348]^x[346]^x[337]^x[332]^x[325]^x[324]^x[321]^x[310]^x[304]^x[299]^x[293]^x[283]^x[282]^x[281]^x[280]^x[273]^x[272]^x[269]^x[262]^x[261]^x[260]^x[254]^x[221]^x[219]^x[217]^x[216]^x[215]^x[212]^x[210]^x[206]^x[205]^x[204]^x[197]^x[193]^x[190]^x[185]^x[184]^x[179]^x[178]^x[175]^x[173]^x[167]^x[164]^x[156]^x[139]^x[135]^x[129]^x[127]^x[126]^x[121]^x[116]^x[115]^x[106]^x[105]^x[97]^x[90]^x[89]^x[79]^x[75]^x[61]^x[59]^x[57]^x[53]^x[52]^x[51]^x[50]^x[47]^x[45]^x[41]^x[39]^x[37]^x[30]^x[25]^x[15]^x[13]^x[9]^x[4]^x[3];
	y[24]=x[379]^x[347]^x[345]^x[336]^x[331]^x[324]^x[323]^x[320]^x[309]^x[303]^x[298]^x[292]^x[282]^x[281]^x[280]^x[279]^x[272]^x[271]^x[268]^x[261]^x[260]^x[259]^x[253]^x[220]^x[218]^x[216]^x[215]^x[214]^x[211]^x[209]^x[205]^x[204]^x[203]^x[196]^x[192]^x[189]^x[184]^x[183]^x[178]^x[177]^x[174]^x[172]^x[166]^x[163]^x[155]^x[138]^x[134]^x[128]^x[127]^x[126]^x[125]^x[120]^x[115]^x[114]^x[106]^x[105]^x[104]^x[96]^x[89]^x[88]^x[78]^x[74]^x[60]^x[58]^x[56]^x[52]^x[51]^x[50]^x[49]^x[46]^x[44]^x[40]^x[38]^x[36]^x[29]^x[24]^x[14]^x[12]^x[8]^x[3]^x[2];
	y[23]=x[378]^x[368]^x[357]^x[346]^x[344]^x[335]^x[323]^x[322]^x[308]^x[302]^x[297]^x[291]^x[281]^x[280]^x[279]^x[278]^x[271]^x[270]^x[267]^x[260]^x[259]^x[258]^x[252]^x[219]^x[217]^x[215]^x[213]^x[210]^x[208]^x[204]^x[202]^x[195]^x[188]^x[183]^x[182]^x[177]^x[176]^x[173]^x[171]^x[165]^x[162]^x[154]^x[137]^x[126]^x[125]^x[124]^x[119]^x[114]^x[113]^x[105]^x[104]^x[103]^x[88]^x[87]^x[77]^x[73]^x[59]^x[57]^x[55]^x[51]^x[50]^x[49]^x[48]^x[45]^x[43]^x[39]^x[37]^x[35]^x[28]^x[23]^x[13]^x[11]^x[7]^x[2]^x[1];
	y[22]=x[377]^x[367]^x[356]^x[345]^x[343]^x[334]^x[322]^x[321]^x[307]^x[301]^x[296]^x[290]^x[280]^x[279]^x[278]^x[277]^x[270]^x[269]^x[266]^x[259]^x[258]^x[257]^x[251]^x[218]^x[216]^x[214]^x[212]^x[209]^x[207]^x[203]^x[201]^x[194]^x[187]^x[182]^x[181]^x[176]^x[175]^x[172]^x[170]^x[164]^x[161]^x[153]^x[136]^x[125]^x[124]^x[123]^x[118]^x[113]^x[112]^x[104]^x[103]^x[102]^x[87]^x[86]^x[76]^x[72]^x[58]^x[56]^x[54]^x[50]^x[49]^x[48]^x[47]^x[44]^x[42]^x[38]^x[36]^x[34]^x[27]^x[22]^x[12]^x[10]^x[6]^x[1]^x[0];
	y[21]=x[376]^x[366]^x[355]^x[344]^x[342]^x[333]^x[321]^x[320]^x[306]^x[300]^x[295]^x[289]^x[279]^x[276]^x[269]^x[268]^x[266]^x[265]^x[258]^x[257]^x[250]^x[217]^x[215]^x[213]^x[211]^x[208]^x[206]^x[203]^x[200]^x[193]^x[192]^x[186]^x[181]^x[180]^x[175]^x[174]^x[171]^x[169]^x[163]^x[160]^x[152]^x[135]^x[124]^x[123]^x[122]^x[117]^x[112]^x[111]^x[103]^x[102]^x[101]^x[86]^x[85]^x[75]^x[71]^x[57]^x[55]^x[53]^x[49]^x[48]^x[47]^x[46]^x[42]^x[41]^x[36]^x[35]^x[33]^x[32]^x[26]^x[21]^x[11]^x[9]^x[5]^x[0];
	y[20]=x[365]^x[354]^x[351]^x[343]^x[341]^x[332]^x[330]^x[320]^x[305]^x[299]^x[294]^x[288]^x[287]^x[286]^x[278]^x[275]^x[268]^x[267]^x[264]^x[257]^x[256]^x[223]^x[222]^x[218]^x[217]^x[214]^x[212]^x[210]^x[206]^x[201]^x[192]^x[191]^x[185]^x[180]^x[179]^x[174]^x[173]^x[168]^x[162]^x[145]^x[134]^x[130]^x[123]^x[122]^x[116]^x[112]^x[110]^x[102]^x[85]^x[84]^x[74]^x[70]^x[63]^x[62]^x[58]^x[56]^x[54]^x[48]^x[46]^x[42]^x[41]^x[40]^x[36]^x[35]^x[34]^x[32]^x[31]^x[20]^x[19]^x[8];
	y[19]=x[351]^x[350]^x[342]^x[340]^x[331]^x[330]^x[329]^x[304]^x[293]^x[287]^x[286]^x[285]^x[277]^x[276]^x[275]^x[274]^x[267]^x[265]^x[263]^x[256]^x[223]^x[221]^x[213]^x[210]^x[209]^x[202]^x[200]^x[199]^x[190]^x[184]^x[179]^x[178]^x[173]^x[172]^x[167]^x[161]^x[144]^x[133]^x[122]^x[115]^x[109]^x[101]^x[84]^x[83]^x[73]^x[69]^x[63]^x[61]^x[57]^x[55]^x[53]^x[51]^x[47]^x[45]^x[42]^x[41]^x[40]^x[39]^x[36]^x[35]^x[34]^x[33]^x[30]^x[19]^x[18]^x[7];
	y[18]=x[350]^x[349]^x[341]^x[339]^x[330]^x[329]^x[328]^x[303]^x[292]^x[287]^x[286]^x[285]^x[284]^x[276]^x[275]^x[274]^x[273]^x[264]^x[262]^x[222]^x[220]^x[212]^x[209]^x[208]^x[201]^x[199]^x[198]^x[189]^x[183]^x[178]^x[177]^x[172]^x[171]^x[166]^x[160]^x[143]^x[132]^x[114]^x[108]^x[83]^x[82]^x[72]^x[68]^x[62]^x[60]^x[56]^x[54]^x[52]^x[50]^x[46]^x[44]^x[41]^x[40]^x[39]^x[38]^x[35]^x[34]^x[33]^x[32]^x[29]^x[18]^x[17]^x[6];
	y[17]=x[349]^x[348]^x[340]^x[338]^x[329]^x[328]^x[327]^x[302]^x[291]^x[286]^x[285]^x[284]^x[283]^x[275]^x[274]^x[273]^x[272]^x[263]^x[261]^x[221]^x[219]^x[214]^x[213]^x[211]^x[202]^x[200]^x[198]^x[196]^x[192]^x[188]^x[182]^x[177]^x[176]^x[171]^x[165]^x[142]^x[131]^x[113]^x[107]^x[82]^x[81]^x[71]^x[67]^x[61]^x[59]^x[55]^x[54]^x[51]^x[49]^x[45]^x[43]^x[42]^x[40]^x[39]^x[38]^x[37]^x[34]^x[33]^x[28]^x[17]^x[16]^x[5];
	y[16]=x[348]^x[347]^x[339]^x[337]^x[328]^x[327]^x[326]^x[301]^x[290]^x[285]^x[284]^x[283]^x[282]^x[274]^x[273]^x[272]^x[271]^x[262]^x[260]^x[220]^x[218]^x[212]^x[210]^x[207]^x[201]^x[199]^x[197]^x[196]^x[195]^x[187]^x[181]^x[176]^x[175]^x[170]^x[164]^x[141]^x[130]^x[112]^x[106]^x[81]^x[80]^x[70]^x[66]^x[60]^x[58]^x[54]^x[50]^x[48]^x[44]^x[42]^x[41]^x[39]^x[38]^x[37]^x[36]^x[33]^x[32]^x[27]^x[16]^x[15]^x[4];
	y[15]=x[347]^x[346]^x[338]^x[336]^x[327]^x[326]^x[325]^x[300]^x[289]^x[284]^x[283]^x[282]^x[281]^x[273]^x[272]^x[271]^x[270]^x[261]^x[259]^x[219]^x[217]^x[213]^x[211]^x[209]^x[207]^x[206]^x[202]^x[200]^x[198]^x[195]^x[194]^x[186]^x[180]^x[175]^x[174]^x[169]^x[163]^x[140]^x[129]^x[111]^x[107]^x[106]^x[105]^x[96]^x[80]^x[79]^x[69]^x[65]^x[59]^x[57]^x[49]^x[47]^x[43]^x[42]^x[41]^x[40]^x[38]^x[37]^x[36]^x[35]^x[32]^x[26]^x[15]^x[14]^x[3];
	y[14]=x[346]^x[345]^x[337]^x[335]^x[326]^x[325]^x[324]^x[299]^x[288]^x[283]^x[282]^x[281]^x[280]^x[272]^x[271]^x[270]^x[269]^x[260]^x[258]^x[218]^x[216]^x[212]^x[210]^x[208]^x[206]^x[205]^x[201]^x[199]^x[197]^x[194]^x[193]^x[185]^x[179]^x[174]^x[173]^x[168]^x[162]^x[139]^x[128]^x[110]^x[105]^x[104]^x[79]^x[78]^x[68]^x[64]^x[58]^x[56]^x[48]^x[46]^x[42]^x[41]^x[40]^x[39]^x[37]^x[36]^x[35]^x[34]^x[25]^x[14]^x[13]^x[2];
	y[13]=x[345]^x[344]^x[336]^x[334]^x[325]^x[324]^x[323]^x[282]^x[281]^x[280]^x[279]^x[271]^x[270]^x[269]^x[268]^x[259]^x[257]^x[217]^x[215]^x[211]^x[209]^x[207]^x[205]^x[204]^x[200]^x[198]^x[196]^x[193]^x[192]^x[184]^x[178]^x[173]^x[172]^x[167]^x[161]^x[109]^x[104]^x[103]^x[78]^x[77]^x[67]^x[57]^x[55]^x[47]^x[45]^x[41]^x[40]^x[39]^x[38]^x[36]^x[35]^x[34]^x[33]^x[24]^x[13]^x[12]^x[1];
	y[12]=x[344]^x[343]^x[335]^x[333]^x[324]^x[323]^x[322]^x[281]^x[280]^x[279]^x[278]^x[270]^x[269]^x[268]^x[267]^x[258]^x[256]^x[216]^x[214]^x[210]^x[208]^x[206]^x[204]^x[199]^x[197]^x[195]^x[183]^x[177]^x[172]^x[171]^x[166]^x[160]^x[108]^x[103]^x[102]^x[77]^x[76]^x[66]^x[56]^x[54]^x[46]^x[44]^x[40]^x[39]^x[38]^x[37]^x[35]^x[34]^x[33]^x[32]^x[23]^x[12]^x[11]^x[0];
	y[11]=x[343]^x[342]^x[334]^x[332]^x[323]^x[322]^x[321]^x[280]^x[279]^x[278]^x[269]^x[267]^x[256]^x[215]^x[214]^x[209]^x[208]^x[205]^x[198]^x[197]^x[194]^x[182]^x[176]^x[171]^x[165]^x[107]^x[102]^x[101]^x[76]^x[75]^x[65]^x[55]^x[54]^x[45]^x[39]^x[38]^x[37]^x[34]^x[33]^x[32]^x[22]^x[11];
	y[10]=x[342]^x[341]^x[333]^x[331]^x[322]^x[321]^x[320]^x[279]^x[278]^x[277]^x[268]^x[267]^x[266]^x[256]^x[214]^x[208]^x[204]^x[202]^x[197]^x[193]^x[181]^x[175]^x[170]^x[164]^x[106]^x[101]^x[100]^x[75]^x[74]^x[64]^x[54]^x[44]^x[42]^x[38]^x[37]^x[36]^x[33]^x[32]^x[21]^x[10];
	y[9]=x[351]^x[341]^x[340]^x[332]^x[321]^x[320]^x[287]^x[286]^x[278]^x[277]^x[275]^x[267]^x[265]^x[221]^x[213]^x[212]^x[211]^x[203]^x[199]^x[192]^x[180]^x[174]^x[169]^x[163]^x[122]^x[105]^x[99]^x[95]^x[73]^x[53]^x[52]^x[51]^x[47]^x[46]^x[45]^x[43]^x[41]^x[37]^x[35]^x[32]^x[20]^x[9];
	y[8]=x[351]^x[350]^x[340]^x[339]^x[331]^x[330]^x[320]^x[285]^x[277]^x[276]^x[275]^x[274]^x[266]^x[264]^x[223]^x[220]^x[212]^x[211]^x[210]^x[198]^x[179]^x[173]^x[168]^x[162]^x[104]^x[98]^x[94]^x[72]^x[63]^x[57]^x[52]^x[50]^x[46]^x[44]^x[40]^x[34]^x[19]^x[8];
	y[7]=x[373]^x[362]^x[351]^x[350]^x[349]^x[339]^x[338]^x[329]^x[284]^x[276]^x[275]^x[274]^x[273]^x[265]^x[263]^x[222]^x[219]^x[211]^x[210]^x[209]^x[197]^x[178]^x[172]^x[167]^x[161]^x[138]^x[132]^x[103]^x[97]^x[93]^x[71]^x[62]^x[56]^x[51]^x[49]^x[45]^x[43]^x[39]^x[33]^x[18]^x[7];
	y[6]=x[372]^x[361]^x[350]^x[349]^x[348]^x[338]^x[337]^x[328]^x[283]^x[275]^x[274]^x[273]^x[272]^x[264]^x[262]^x[221]^x[218]^x[210]^x[209]^x[208]^x[196]^x[177]^x[171]^x[166]^x[160]^x[137]^x[131]^x[102]^x[96]^x[92]^x[70]^x[61]^x[55]^x[50]^x[48]^x[44]^x[42]^x[38]^x[32]^x[17]^x[6];
	y[5]=x[371]^x[360]^x[349]^x[348]^x[347]^x[337]^x[336]^x[327]^x[282]^x[274]^x[273]^x[271]^x[263]^x[245]^x[234]^x[220]^x[217]^x[214]^x[209]^x[207]^x[197]^x[195]^x[192]^x[176]^x[165]^x[136]^x[130]^x[118]^x[108]^x[107]^x[106]^x[101]^x[97]^x[96]^x[91]^x[69]^x[60]^x[49]^x[47]^x[43]^x[41]^x[32]^x[16]^x[10]^x[5]^x[4];
	y[4]=x[370]^x[359]^x[348]^x[347]^x[346]^x[336]^x[335]^x[326]^x[281]^x[273]^x[272]^x[271]^x[270]^x[262]^x[260]^x[244]^x[233]^x[219]^x[216]^x[213]^x[208]^x[206]^x[202]^x[196]^x[194]^x[175]^x[164]^x[135]^x[129]^x[107]^x[106]^x[105]^x[100]^x[96]^x[90]^x[68]^x[59]^x[48]^x[46]^x[40]^x[36]^x[15]^x[9]^x[4]^x[3];
	y[3]=x[369]^x[358]^x[347]^x[346]^x[345]^x[335]^x[334]^x[325]^x[280]^x[272]^x[271]^x[270]^x[269]^x[261]^x[259]^x[243]^x[232]^x[218]^x[215]^x[212]^x[207]^x[205]^x[201]^x[195]^x[193]^x[174]^x[163]^x[134]^x[128]^x[106]^x[105]^x[104]^x[99]^x[89]^x[67]^x[58]^x[47]^x[45]^x[39]^x[35]^x[14]^x[8]^x[3]^x[2];
	y[2]=x[368]^x[357]^x[346]^x[345]^x[344]^x[334]^x[333]^x[324]^x[279]^x[271]^x[270]^x[269]^x[268]^x[260]^x[258]^x[242]^x[231]^x[217]^x[214]^x[211]^x[206]^x[204]^x[200]^x[194]^x[192]^x[173]^x[162]^x[133]^x[105]^x[104]^x[103]^x[98]^x[88]^x[66]^x[57]^x[46]^x[44]^x[38]^x[34]^x[13]^x[7]^x[2]^x[1];
	y[1]=x[345]^x[344]^x[343]^x[333]^x[332]^x[323]^x[278]^x[270]^x[269]^x[268]^x[267]^x[259]^x[257]^x[241]^x[230]^x[216]^x[210]^x[205]^x[203]^x[199]^x[193]^x[172]^x[161]^x[104]^x[103]^x[102]^x[97]^x[87]^x[65]^x[56]^x[45]^x[43]^x[37]^x[33]^x[12]^x[6]^x[1]^x[0];
	y[0]=x[344]^x[343]^x[342]^x[332]^x[331]^x[322]^x[278]^x[269]^x[268]^x[267]^x[258]^x[240]^x[229]^x[215]^x[209]^x[204]^x[203]^x[198]^x[171]^x[160]^x[103]^x[102]^x[101]^x[96]^x[86]^x[64]^x[55]^x[44]^x[43]^x[37]^x[11]^x[5]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint62(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[373]^x[372]^x[371]^x[363]^x[361]^x[352]^x[333]^x[322]^x[311]^x[306]^x[301]^x[298]^x[295]^x[290]^x[288]^x[284]^x[278]^x[273]^x[267]^x[255]^x[254]^x[247]^x[246]^x[245]^x[244]^x[243]^x[235]^x[225]^x[186]^x[185]^x[181]^x[176]^x[174]^x[172]^x[171]^x[170]^x[167]^x[165]^x[161]^x[124]^x[113]^x[98]^x[95]^x[91]^x[90]^x[89]^x[80]^x[71]^x[70]^x[65]^x[63]^x[53]^x[49]^x[43]^x[37]^x[32]^x[26]^x[25]^x[21]^x[20]^x[19]^x[16]^x[15]^x[13]^x[12]^x[11]^x[6]^x[1]^x[0];
	y[30]=x[383]^x[382]^x[372]^x[371]^x[370]^x[360]^x[319]^x[310]^x[305]^x[300]^x[298]^x[297]^x[294]^x[289]^x[283]^x[277]^x[272]^x[266]^x[254]^x[253]^x[246]^x[245]^x[244]^x[242]^x[234]^x[233]^x[224]^x[190]^x[189]^x[178]^x[171]^x[170]^x[166]^x[160]^x[123]^x[112]^x[94]^x[88]^x[70]^x[69]^x[64]^x[63]^x[62]^x[52]^x[48]^x[36]^x[30]^x[24]^x[18]^x[12]^x[11]^x[10]^x[5]^x[4]^x[0];
	y[29]=x[382]^x[381]^x[371]^x[370]^x[369]^x[359]^x[342]^x[320]^x[318]^x[309]^x[304]^x[299]^x[297]^x[296]^x[293]^x[288]^x[282]^x[276]^x[271]^x[265]^x[255]^x[254]^x[253]^x[252]^x[245]^x[244]^x[241]^x[234]^x[233]^x[232]^x[191]^x[189]^x[188]^x[177]^x[169]^x[165]^x[122]^x[111]^x[107]^x[101]^x[96]^x[93]^x[87]^x[69]^x[62]^x[61]^x[51]^x[47]^x[35]^x[31]^x[29]^x[25]^x[23]^x[19]^x[17]^x[13]^x[11]^x[9]^x[3];
	y[28]=x[381]^x[380]^x[370]^x[369]^x[368]^x[358]^x[341]^x[330]^x[319]^x[317]^x[308]^x[303]^x[296]^x[295]^x[292]^x[281]^x[275]^x[270]^x[264]^x[254]^x[253]^x[252]^x[251]^x[244]^x[243]^x[240]^x[233]^x[232]^x[231]^x[190]^x[188]^x[187]^x[176]^x[168]^x[164]^x[121]^x[110]^x[106]^x[100]^x[92]^x[86]^x[68]^x[61]^x[60]^x[50]^x[46]^x[34]^x[30]^x[28]^x[24]^x[22]^x[18]^x[16]^x[12]^x[10]^x[8]^x[2];
	y[27]=x[380]^x[379]^x[369]^x[368]^x[367]^x[357]^x[340]^x[329]^x[318]^x[316]^x[307]^x[302]^x[295]^x[294]^x[291]^x[280]^x[274]^x[269]^x[263]^x[253]^x[252]^x[251]^x[250]^x[243]^x[242]^x[239]^x[232]^x[231]^x[230]^x[189]^x[187]^x[186]^x[175]^x[167]^x[163]^x[120]^x[109]^x[105]^x[99]^x[91]^x[85]^x[67]^x[60]^x[59]^x[49]^x[45]^x[33]^x[29]^x[27]^x[23]^x[21]^x[17]^x[15]^x[11]^x[9]^x[7]^x[1];
	y[26]=x[383]^x[379]^x[378]^x[377]^x[368]^x[367]^x[366]^x[356]^x[349]^x[339]^x[328]^x[317]^x[315]^x[306]^x[301]^x[294]^x[293]^x[290]^x[279]^x[273]^x[268]^x[262]^x[252]^x[251]^x[249]^x[242]^x[241]^x[238]^x[231]^x[230]^x[229]^x[223]^x[191]^x[190]^x[188]^x[184]^x[181]^x[180]^x[179]^x[175]^x[173]^x[171]^x[166]^x[162]^x[160]^x[147]^x[125]^x[108]^x[95]^x[90]^x[86]^x[85]^x[84]^x[75]^x[74]^x[66]^x[59]^x[58]^x[48]^x[44]^x[32]^x[31]^x[30]^x[28]^x[22]^x[21]^x[20]^x[19]^x[16]^x[14]^x[11]^x[10]^x[8]^x[6]^x[5];
	y[25]=x[382]^x[378]^x[377]^x[376]^x[367]^x[366]^x[365]^x[355]^x[348]^x[316]^x[314]^x[305]^x[300]^x[293]^x[292]^x[289]^x[278]^x[272]^x[267]^x[261]^x[251]^x[250]^x[249]^x[248]^x[241]^x[240]^x[237]^x[230]^x[229]^x[228]^x[222]^x[189]^x[187]^x[185]^x[184]^x[183]^x[180]^x[178]^x[174]^x[173]^x[172]^x[165]^x[161]^x[146]^x[124]^x[107]^x[103]^x[97]^x[95]^x[94]^x[89]^x[84]^x[83]^x[74]^x[73]^x[65]^x[58]^x[57]^x[47]^x[43]^x[29]^x[27]^x[25]^x[21]^x[20]^x[19]^x[18]^x[15]^x[13]^x[9]^x[7]^x[5];
	y[24]=x[381]^x[377]^x[376]^x[375]^x[366]^x[365]^x[364]^x[354]^x[347]^x[315]^x[313]^x[304]^x[299]^x[292]^x[291]^x[288]^x[277]^x[271]^x[266]^x[260]^x[250]^x[249]^x[248]^x[247]^x[240]^x[239]^x[236]^x[229]^x[228]^x[227]^x[221]^x[188]^x[186]^x[184]^x[183]^x[182]^x[179]^x[177]^x[173]^x[172]^x[171]^x[164]^x[160]^x[145]^x[123]^x[106]^x[102]^x[96]^x[95]^x[94]^x[93]^x[88]^x[83]^x[82]^x[74]^x[73]^x[72]^x[64]^x[57]^x[56]^x[46]^x[42]^x[28]^x[26]^x[24]^x[20]^x[19]^x[18]^x[17]^x[14]^x[12]^x[8]^x[6]^x[4];
	y[23]=x[380]^x[376]^x[375]^x[374]^x[365]^x[364]^x[363]^x[353]^x[346]^x[336]^x[325]^x[314]^x[312]^x[303]^x[291]^x[290]^x[276]^x[270]^x[265]^x[259]^x[249]^x[248]^x[247]^x[246]^x[239]^x[238]^x[235]^x[228]^x[227]^x[226]^x[220]^x[187]^x[185]^x[183]^x[181]^x[178]^x[176]^x[172]^x[170]^x[163]^x[144]^x[122]^x[105]^x[94]^x[93]^x[92]^x[87]^x[82]^x[81]^x[73]^x[72]^x[71]^x[56]^x[55]^x[45]^x[41]^x[27]^x[25]^x[23]^x[19]^x[18]^x[17]^x[16]^x[13]^x[11]^x[7]^x[5]^x[3];
	y[22]=x[379]^x[375]^x[374]^x[373]^x[364]^x[363]^x[362]^x[352]^x[345]^x[335]^x[324]^x[313]^x[311]^x[302]^x[290]^x[289]^x[275]^x[269]^x[264]^x[258]^x[248]^x[247]^x[246]^x[245]^x[238]^x[237]^x[234]^x[227]^x[226]^x[225]^x[219]^x[186]^x[184]^x[182]^x[180]^x[177]^x[175]^x[171]^x[169]^x[162]^x[143]^x[121]^x[104]^x[93]^x[92]^x[91]^x[86]^x[81]^x[80]^x[72]^x[71]^x[70]^x[55]^x[54]^x[44]^x[40]^x[26]^x[24]^x[22]^x[18]^x[17]^x[16]^x[15]^x[12]^x[10]^x[6]^x[4]^x[2];
	y[21]=x[378]^x[374]^x[373]^x[372]^x[363]^x[361]^x[344]^x[334]^x[323]^x[312]^x[310]^x[301]^x[289]^x[288]^x[274]^x[268]^x[263]^x[257]^x[247]^x[244]^x[237]^x[236]^x[234]^x[233]^x[226]^x[225]^x[218]^x[185]^x[183]^x[181]^x[179]^x[176]^x[174]^x[171]^x[168]^x[161]^x[160]^x[142]^x[120]^x[103]^x[92]^x[91]^x[90]^x[85]^x[80]^x[79]^x[71]^x[70]^x[69]^x[54]^x[53]^x[43]^x[39]^x[25]^x[23]^x[21]^x[17]^x[16]^x[15]^x[14]^x[10]^x[9]^x[4]^x[3]^x[1]^x[0];
	y[20]=x[382]^x[373]^x[372]^x[362]^x[360]^x[333]^x[322]^x[319]^x[311]^x[309]^x[300]^x[298]^x[288]^x[273]^x[267]^x[262]^x[256]^x[255]^x[254]^x[246]^x[243]^x[236]^x[235]^x[232]^x[225]^x[224]^x[191]^x[190]^x[186]^x[185]^x[182]^x[180]^x[178]^x[174]^x[169]^x[160]^x[113]^x[102]^x[98]^x[91]^x[90]^x[84]^x[80]^x[78]^x[70]^x[53]^x[52]^x[42]^x[38]^x[31]^x[30]^x[26]^x[24]^x[22]^x[16]^x[14]^x[10]^x[9]^x[8]^x[4]^x[3]^x[2]^x[0];
	y[19]=x[381]^x[372]^x[371]^x[361]^x[359]^x[319]^x[318]^x[310]^x[308]^x[299]^x[298]^x[297]^x[272]^x[261]^x[255]^x[254]^x[253]^x[245]^x[244]^x[243]^x[242]^x[235]^x[233]^x[231]^x[224]^x[191]^x[189]^x[181]^x[178]^x[177]^x[170]^x[168]^x[167]^x[112]^x[101]^x[90]^x[83]^x[77]^x[69]^x[52]^x[51]^x[41]^x[37]^x[31]^x[29]^x[25]^x[23]^x[21]^x[19]^x[15]^x[13]^x[10]^x[9]^x[8]^x[7]^x[4]^x[3]^x[2]^x[1];
	y[18]=x[380]^x[371]^x[370]^x[360]^x[358]^x[318]^x[317]^x[309]^x[307]^x[298]^x[297]^x[296]^x[271]^x[260]^x[255]^x[254]^x[253]^x[252]^x[244]^x[243]^x[242]^x[241]^x[232]^x[230]^x[190]^x[188]^x[180]^x[177]^x[176]^x[169]^x[167]^x[166]^x[111]^x[100]^x[82]^x[76]^x[51]^x[50]^x[40]^x[36]^x[30]^x[28]^x[24]^x[22]^x[20]^x[18]^x[14]^x[12]^x[9]^x[8]^x[7]^x[6]^x[3]^x[2]^x[1]^x[0];
	y[17]=x[379]^x[370]^x[369]^x[359]^x[357]^x[317]^x[316]^x[308]^x[306]^x[297]^x[296]^x[295]^x[270]^x[259]^x[254]^x[253]^x[252]^x[251]^x[243]^x[242]^x[241]^x[240]^x[231]^x[229]^x[189]^x[187]^x[182]^x[181]^x[179]^x[170]^x[168]^x[166]^x[164]^x[160]^x[138]^x[110]^x[99]^x[81]^x[75]^x[50]^x[49]^x[39]^x[35]^x[29]^x[27]^x[23]^x[22]^x[19]^x[17]^x[13]^x[11]^x[10]^x[8]^x[7]^x[6]^x[5]^x[2]^x[1];
	y[16]=x[378]^x[369]^x[368]^x[358]^x[356]^x[316]^x[315]^x[307]^x[305]^x[296]^x[295]^x[294]^x[269]^x[258]^x[253]^x[252]^x[251]^x[250]^x[242]^x[241]^x[240]^x[239]^x[230]^x[228]^x[188]^x[186]^x[180]^x[178]^x[175]^x[169]^x[167]^x[165]^x[164]^x[163]^x[137]^x[109]^x[98]^x[80]^x[74]^x[49]^x[48]^x[38]^x[34]^x[28]^x[26]^x[22]^x[18]^x[16]^x[12]^x[10]^x[9]^x[7]^x[6]^x[5]^x[4]^x[1]^x[0];
	y[15]=x[377]^x[368]^x[367]^x[357]^x[355]^x[315]^x[314]^x[306]^x[304]^x[295]^x[294]^x[293]^x[268]^x[257]^x[252]^x[251]^x[250]^x[249]^x[241]^x[240]^x[239]^x[238]^x[229]^x[227]^x[187]^x[185]^x[181]^x[179]^x[177]^x[175]^x[174]^x[170]^x[168]^x[166]^x[163]^x[162]^x[136]^x[108]^x[97]^x[79]^x[75]^x[74]^x[73]^x[64]^x[48]^x[47]^x[37]^x[33]^x[27]^x[25]^x[17]^x[15]^x[11]^x[10]^x[9]^x[8]^x[6]^x[5]^x[4]^x[3]^x[0];
	y[14]=x[376]^x[367]^x[366]^x[356]^x[354]^x[314]^x[313]^x[305]^x[303]^x[294]^x[293]^x[292]^x[267]^x[256]^x[251]^x[250]^x[249]^x[248]^x[240]^x[239]^x[238]^x[237]^x[228]^x[226]^x[186]^x[184]^x[180]^x[178]^x[176]^x[174]^x[173]^x[169]^x[167]^x[165]^x[162]^x[161]^x[135]^x[107]^x[96]^x[78]^x[73]^x[72]^x[47]^x[46]^x[36]^x[32]^x[26]^x[24]^x[16]^x[14]^x[10]^x[9]^x[8]^x[7]^x[5]^x[4]^x[3]^x[2];
	y[13]=x[375]^x[366]^x[365]^x[355]^x[353]^x[313]^x[312]^x[304]^x[302]^x[293]^x[292]^x[291]^x[250]^x[249]^x[248]^x[247]^x[239]^x[238]^x[237]^x[236]^x[227]^x[225]^x[185]^x[183]^x[179]^x[177]^x[175]^x[173]^x[172]^x[168]^x[166]^x[164]^x[161]^x[160]^x[134]^x[77]^x[72]^x[71]^x[46]^x[45]^x[35]^x[25]^x[23]^x[15]^x[13]^x[9]^x[8]^x[7]^x[6]^x[4]^x[3]^x[2]^x[1];
	y[12]=x[374]^x[365]^x[364]^x[354]^x[352]^x[312]^x[311]^x[303]^x[301]^x[292]^x[291]^x[290]^x[249]^x[248]^x[247]^x[246]^x[238]^x[237]^x[236]^x[235]^x[226]^x[224]^x[184]^x[182]^x[178]^x[176]^x[174]^x[172]^x[167]^x[165]^x[163]^x[133]^x[76]^x[71]^x[70]^x[45]^x[44]^x[34]^x[24]^x[22]^x[14]^x[12]^x[8]^x[7]^x[6]^x[5]^x[3]^x[2]^x[1]^x[0];
	y[11]=x[364]^x[363]^x[353]^x[311]^x[310]^x[302]^x[300]^x[291]^x[290]^x[289]^x[248]^x[247]^x[246]^x[237]^x[235]^x[224]^x[183]^x[182]^x[177]^x[176]^x[173]^x[166]^x[165]^x[162]^x[75]^x[70]^x[69]^x[44]^x[43]^x[33]^x[23]^x[22]^x[13]^x[7]^x[6]^x[5]^x[2]^x[1]^x[0];
	y[10]=x[363]^x[362]^x[352]^x[310]^x[309]^x[301]^x[299]^x[290]^x[289]^x[288]^x[247]^x[246]^x[245]^x[236]^x[235]^x[234]^x[224]^x[182]^x[176]^x[172]^x[170]^x[165]^x[161]^x[74]^x[69]^x[68]^x[43]^x[42]^x[32]^x[22]^x[12]^x[10]^x[6]^x[5]^x[4]^x[1]^x[0];
	y[9]=x[383]^x[361]^x[319]^x[309]^x[308]^x[300]^x[289]^x[288]^x[255]^x[254]^x[246]^x[245]^x[243]^x[235]^x[233]^x[189]^x[181]^x[180]^x[179]^x[171]^x[167]^x[160]^x[90]^x[73]^x[67]^x[63]^x[41]^x[21]^x[20]^x[19]^x[15]^x[14]^x[13]^x[11]^x[9]^x[5]^x[3]^x[0];
	y[8]=x[382]^x[360]^x[319]^x[318]^x[308]^x[307]^x[299]^x[298]^x[288]^x[253]^x[245]^x[244]^x[243]^x[242]^x[234]^x[232]^x[191]^x[188]^x[180]^x[179]^x[178]^x[166]^x[72]^x[66]^x[62]^x[40]^x[31]^x[25]^x[20]^x[18]^x[14]^x[12]^x[8]^x[2];
	y[7]=x[381]^x[359]^x[341]^x[330]^x[319]^x[318]^x[317]^x[307]^x[306]^x[297]^x[252]^x[244]^x[243]^x[242]^x[241]^x[233]^x[231]^x[190]^x[187]^x[179]^x[178]^x[177]^x[165]^x[106]^x[100]^x[71]^x[65]^x[61]^x[39]^x[30]^x[24]^x[19]^x[17]^x[13]^x[11]^x[7]^x[1];
	y[6]=x[380]^x[358]^x[340]^x[329]^x[318]^x[317]^x[316]^x[306]^x[305]^x[296]^x[251]^x[243]^x[242]^x[241]^x[240]^x[232]^x[230]^x[189]^x[186]^x[178]^x[177]^x[176]^x[164]^x[105]^x[99]^x[70]^x[64]^x[60]^x[38]^x[29]^x[23]^x[18]^x[16]^x[12]^x[10]^x[6]^x[0];
	y[5]=x[379]^x[373]^x[367]^x[362]^x[357]^x[356]^x[339]^x[328]^x[317]^x[316]^x[315]^x[305]^x[304]^x[295]^x[250]^x[242]^x[241]^x[239]^x[231]^x[213]^x[202]^x[188]^x[185]^x[182]^x[177]^x[175]^x[165]^x[163]^x[160]^x[104]^x[98]^x[86]^x[76]^x[75]^x[74]^x[69]^x[65]^x[64]^x[59]^x[37]^x[28]^x[17]^x[15]^x[11]^x[9]^x[0];
	y[4]=x[378]^x[372]^x[366]^x[361]^x[356]^x[355]^x[338]^x[327]^x[316]^x[315]^x[314]^x[304]^x[303]^x[294]^x[249]^x[241]^x[240]^x[239]^x[238]^x[230]^x[228]^x[212]^x[201]^x[187]^x[184]^x[181]^x[176]^x[174]^x[170]^x[164]^x[162]^x[103]^x[97]^x[75]^x[74]^x[73]^x[68]^x[64]^x[58]^x[36]^x[27]^x[16]^x[14]^x[8]^x[4];
	y[3]=x[377]^x[371]^x[365]^x[360]^x[355]^x[354]^x[337]^x[326]^x[315]^x[314]^x[313]^x[303]^x[302]^x[293]^x[248]^x[240]^x[239]^x[238]^x[237]^x[229]^x[227]^x[211]^x[200]^x[186]^x[183]^x[180]^x[175]^x[173]^x[169]^x[163]^x[161]^x[102]^x[96]^x[74]^x[73]^x[72]^x[67]^x[57]^x[35]^x[26]^x[15]^x[13]^x[7]^x[3];
	y[2]=x[376]^x[370]^x[364]^x[359]^x[354]^x[353]^x[336]^x[325]^x[314]^x[313]^x[312]^x[302]^x[301]^x[292]^x[247]^x[239]^x[238]^x[237]^x[236]^x[228]^x[226]^x[210]^x[199]^x[185]^x[182]^x[179]^x[174]^x[172]^x[168]^x[162]^x[160]^x[101]^x[73]^x[72]^x[71]^x[66]^x[56]^x[34]^x[25]^x[14]^x[12]^x[6]^x[2];
	y[1]=x[375]^x[369]^x[363]^x[358]^x[353]^x[352]^x[313]^x[312]^x[311]^x[301]^x[300]^x[291]^x[246]^x[238]^x[237]^x[236]^x[235]^x[227]^x[225]^x[209]^x[198]^x[184]^x[178]^x[173]^x[171]^x[167]^x[161]^x[72]^x[71]^x[70]^x[65]^x[55]^x[33]^x[24]^x[13]^x[11]^x[5]^x[1];
	y[0]=x[374]^x[368]^x[357]^x[352]^x[312]^x[311]^x[310]^x[300]^x[299]^x[290]^x[246]^x[237]^x[236]^x[235]^x[226]^x[208]^x[197]^x[183]^x[177]^x[172]^x[171]^x[166]^x[71]^x[70]^x[69]^x[64]^x[54]^x[32]^x[23]^x[12]^x[11]^x[5];
	return y;
endfunction

(* noinline *)
function Bit#(32) randint63(Bit#(384) x);
	Bit#(32) y = 0;
	y[31]=x[383]^x[382]^x[379]^x[377]^x[376]^x[375]^x[374]^x[373]^x[372]^x[371]^x[369]^x[365]^x[363]^x[358]^x[357]^x[356]^x[353]^x[351]^x[341]^x[340]^x[339]^x[331]^x[329]^x[320]^x[301]^x[290]^x[279]^x[274]^x[269]^x[266]^x[263]^x[258]^x[256]^x[252]^x[246]^x[241]^x[235]^x[223]^x[222]^x[215]^x[214]^x[213]^x[212]^x[211]^x[203]^x[193]^x[137]^x[92]^x[81]^x[66]^x[63]^x[59]^x[58]^x[57]^x[48]^x[39]^x[38]^x[33]^x[31]^x[21]^x[17]^x[11]^x[5]^x[0];
	y[30]=x[382]^x[381]^x[376]^x[375]^x[374]^x[373]^x[372]^x[370]^x[368]^x[367]^x[366]^x[364]^x[362]^x[361]^x[357]^x[356]^x[355]^x[352]^x[351]^x[350]^x[340]^x[339]^x[338]^x[328]^x[287]^x[278]^x[273]^x[268]^x[266]^x[265]^x[262]^x[257]^x[251]^x[245]^x[240]^x[234]^x[222]^x[221]^x[214]^x[213]^x[212]^x[210]^x[202]^x[201]^x[192]^x[157]^x[146]^x[91]^x[80]^x[62]^x[56]^x[38]^x[37]^x[32]^x[31]^x[30]^x[20]^x[16]^x[4];
	y[29]=x[383]^x[382]^x[381]^x[380]^x[377]^x[376]^x[375]^x[374]^x[373]^x[372]^x[369]^x[367]^x[366]^x[363]^x[362]^x[361]^x[360]^x[356]^x[355]^x[354]^x[350]^x[349]^x[339]^x[338]^x[337]^x[327]^x[310]^x[288]^x[286]^x[277]^x[272]^x[267]^x[265]^x[264]^x[261]^x[256]^x[250]^x[244]^x[239]^x[233]^x[223]^x[222]^x[221]^x[220]^x[213]^x[212]^x[209]^x[202]^x[201]^x[200]^x[156]^x[145]^x[135]^x[90]^x[79]^x[75]^x[69]^x[64]^x[61]^x[55]^x[37]^x[30]^x[29]^x[19]^x[15]^x[3];
	y[28]=x[382]^x[381]^x[380]^x[379]^x[376]^x[375]^x[374]^x[373]^x[372]^x[371]^x[368]^x[366]^x[365]^x[362]^x[361]^x[360]^x[359]^x[355]^x[354]^x[353]^x[349]^x[348]^x[338]^x[337]^x[336]^x[326]^x[309]^x[298]^x[287]^x[285]^x[276]^x[271]^x[264]^x[263]^x[260]^x[249]^x[243]^x[238]^x[232]^x[222]^x[221]^x[220]^x[219]^x[212]^x[211]^x[208]^x[201]^x[200]^x[199]^x[155]^x[144]^x[134]^x[89]^x[78]^x[74]^x[68]^x[60]^x[54]^x[36]^x[29]^x[28]^x[18]^x[14]^x[2];
	y[27]=x[381]^x[380]^x[379]^x[378]^x[375]^x[374]^x[373]^x[372]^x[371]^x[370]^x[367]^x[365]^x[364]^x[361]^x[360]^x[359]^x[358]^x[354]^x[353]^x[352]^x[348]^x[347]^x[337]^x[336]^x[335]^x[325]^x[308]^x[297]^x[286]^x[284]^x[275]^x[270]^x[263]^x[262]^x[259]^x[248]^x[242]^x[237]^x[231]^x[221]^x[220]^x[219]^x[218]^x[211]^x[210]^x[207]^x[200]^x[199]^x[198]^x[154]^x[143]^x[133]^x[88]^x[77]^x[73]^x[67]^x[59]^x[53]^x[35]^x[28]^x[27]^x[17]^x[13]^x[1];
	y[26]=x[380]^x[379]^x[377]^x[373]^x[370]^x[369]^x[366]^x[364]^x[361]^x[360]^x[359]^x[358]^x[357]^x[353]^x[352]^x[351]^x[347]^x[346]^x[345]^x[336]^x[335]^x[334]^x[324]^x[317]^x[307]^x[296]^x[285]^x[283]^x[274]^x[269]^x[262]^x[261]^x[258]^x[247]^x[241]^x[236]^x[230]^x[220]^x[219]^x[217]^x[210]^x[209]^x[206]^x[199]^x[198]^x[197]^x[191]^x[153]^x[132]^x[115]^x[93]^x[76]^x[63]^x[58]^x[54]^x[53]^x[52]^x[43]^x[42]^x[34]^x[27]^x[26]^x[16]^x[12]^x[0];
	y[25]=x[383]^x[382]^x[379]^x[378]^x[377]^x[376]^x[373]^x[369]^x[368]^x[365]^x[363]^x[361]^x[360]^x[359]^x[358]^x[357]^x[356]^x[352]^x[350]^x[346]^x[345]^x[344]^x[335]^x[334]^x[333]^x[323]^x[316]^x[284]^x[282]^x[273]^x[268]^x[261]^x[260]^x[257]^x[246]^x[240]^x[235]^x[229]^x[219]^x[218]^x[217]^x[216]^x[209]^x[208]^x[205]^x[198]^x[197]^x[196]^x[190]^x[152]^x[141]^x[131]^x[114]^x[92]^x[75]^x[71]^x[65]^x[63]^x[62]^x[57]^x[52]^x[51]^x[42]^x[41]^x[33]^x[26]^x[25]^x[15]^x[11];
	y[24]=x[383]^x[382]^x[381]^x[378]^x[377]^x[376]^x[375]^x[372]^x[368]^x[367]^x[364]^x[360]^x[359]^x[358]^x[357]^x[356]^x[355]^x[349]^x[345]^x[344]^x[343]^x[334]^x[333]^x[332]^x[322]^x[315]^x[283]^x[281]^x[272]^x[267]^x[260]^x[259]^x[256]^x[245]^x[239]^x[234]^x[228]^x[218]^x[217]^x[216]^x[215]^x[208]^x[207]^x[204]^x[197]^x[196]^x[195]^x[189]^x[151]^x[140]^x[130]^x[113]^x[91]^x[74]^x[70]^x[64]^x[63]^x[62]^x[61]^x[56]^x[51]^x[50]^x[42]^x[41]^x[40]^x[32]^x[25]^x[24]^x[14]^x[10];
	y[23]=x[382]^x[381]^x[380]^x[377]^x[376]^x[375]^x[374]^x[371]^x[367]^x[366]^x[363]^x[359]^x[358]^x[357]^x[356]^x[355]^x[354]^x[348]^x[344]^x[343]^x[342]^x[333]^x[332]^x[331]^x[321]^x[314]^x[304]^x[293]^x[282]^x[280]^x[271]^x[259]^x[258]^x[244]^x[238]^x[233]^x[227]^x[217]^x[216]^x[215]^x[214]^x[207]^x[206]^x[203]^x[196]^x[195]^x[194]^x[188]^x[129]^x[112]^x[90]^x[73]^x[62]^x[61]^x[60]^x[55]^x[50]^x[49]^x[41]^x[40]^x[39]^x[24]^x[23]^x[13]^x[9];
	y[22]=x[381]^x[380]^x[379]^x[376]^x[375]^x[374]^x[373]^x[370]^x[366]^x[365]^x[362]^x[358]^x[357]^x[356]^x[355]^x[354]^x[353]^x[347]^x[343]^x[342]^x[341]^x[332]^x[331]^x[330]^x[320]^x[313]^x[303]^x[292]^x[281]^x[279]^x[270]^x[258]^x[257]^x[243]^x[237]^x[232]^x[226]^x[216]^x[215]^x[214]^x[213]^x[206]^x[205]^x[202]^x[195]^x[194]^x[193]^x[187]^x[128]^x[111]^x[89]^x[72]^x[61]^x[60]^x[59]^x[54]^x[49]^x[48]^x[40]^x[39]^x[38]^x[23]^x[22]^x[12]^x[8];
	y[21]=x[380]^x[379]^x[378]^x[375]^x[372]^x[369]^x[368]^x[367]^x[365]^x[364]^x[362]^x[361]^x[355]^x[354]^x[353]^x[346]^x[342]^x[341]^x[340]^x[331]^x[329]^x[312]^x[302]^x[291]^x[280]^x[278]^x[269]^x[257]^x[256]^x[242]^x[236]^x[231]^x[225]^x[215]^x[212]^x[205]^x[204]^x[202]^x[201]^x[194]^x[193]^x[186]^x[110]^x[88]^x[71]^x[60]^x[59]^x[58]^x[53]^x[48]^x[47]^x[39]^x[38]^x[37]^x[22]^x[21]^x[11]^x[7];
	y[20]=x[383]^x[382]^x[379]^x[378]^x[377]^x[376]^x[374]^x[371]^x[367]^x[366]^x[365]^x[364]^x[363]^x[360]^x[357]^x[356]^x[354]^x[353]^x[352]^x[350]^x[341]^x[340]^x[330]^x[328]^x[301]^x[290]^x[287]^x[279]^x[277]^x[268]^x[266]^x[256]^x[241]^x[235]^x[230]^x[224]^x[223]^x[222]^x[214]^x[211]^x[204]^x[203]^x[200]^x[193]^x[192]^x[81]^x[70]^x[66]^x[59]^x[58]^x[52]^x[48]^x[46]^x[38]^x[21]^x[20]^x[10]^x[6];
	y[19]=x[383]^x[382]^x[381]^x[378]^x[377]^x[376]^x[375]^x[373]^x[372]^x[371]^x[370]^x[367]^x[366]^x[365]^x[364]^x[363]^x[361]^x[359]^x[355]^x[353]^x[352]^x[349]^x[340]^x[339]^x[329]^x[327]^x[287]^x[286]^x[278]^x[276]^x[267]^x[266]^x[265]^x[240]^x[229]^x[223]^x[222]^x[221]^x[213]^x[212]^x[211]^x[210]^x[203]^x[201]^x[199]^x[192]^x[146]^x[135]^x[80]^x[69]^x[58]^x[51]^x[45]^x[37]^x[20]^x[19]^x[9]^x[5];
	y[18]=x[383]^x[382]^x[381]^x[380]^x[377]^x[376]^x[375]^x[374]^x[372]^x[371]^x[370]^x[369]^x[366]^x[365]^x[364]^x[363]^x[360]^x[358]^x[354]^x[352]^x[348]^x[339]^x[338]^x[328]^x[326]^x[286]^x[285]^x[277]^x[275]^x[266]^x[265]^x[264]^x[239]^x[228]^x[223]^x[222]^x[221]^x[220]^x[212]^x[211]^x[210]^x[209]^x[200]^x[198]^x[145]^x[134]^x[79]^x[68]^x[50]^x[44]^x[19]^x[18]^x[8]^x[4];
	y[17]=x[382]^x[381]^x[380]^x[379]^x[376]^x[375]^x[373]^x[371]^x[370]^x[369]^x[368]^x[365]^x[363]^x[362]^x[359]^x[357]^x[347]^x[338]^x[337]^x[327]^x[325]^x[285]^x[284]^x[276]^x[274]^x[265]^x[264]^x[263]^x[238]^x[227]^x[222]^x[221]^x[220]^x[219]^x[211]^x[210]^x[209]^x[208]^x[199]^x[197]^x[144]^x[106]^x[78]^x[67]^x[49]^x[43]^x[18]^x[17]^x[7]^x[3];
	y[16]=x[381]^x[380]^x[379]^x[378]^x[375]^x[374]^x[373]^x[372]^x[370]^x[369]^x[368]^x[367]^x[364]^x[363]^x[362]^x[361]^x[358]^x[356]^x[352]^x[346]^x[337]^x[336]^x[326]^x[324]^x[284]^x[283]^x[275]^x[273]^x[264]^x[263]^x[262]^x[237]^x[226]^x[221]^x[220]^x[219]^x[218]^x[210]^x[209]^x[208]^x[207]^x[198]^x[196]^x[143]^x[132]^x[105]^x[77]^x[66]^x[48]^x[42]^x[17]^x[16]^x[6]^x[2];
	y[15]=x[380]^x[379]^x[378]^x[377]^x[374]^x[373]^x[372]^x[371]^x[369]^x[368]^x[367]^x[366]^x[362]^x[361]^x[360]^x[357]^x[355]^x[352]^x[345]^x[336]^x[335]^x[325]^x[323]^x[283]^x[282]^x[274]^x[272]^x[263]^x[262]^x[261]^x[236]^x[225]^x[220]^x[219]^x[218]^x[217]^x[209]^x[208]^x[207]^x[206]^x[197]^x[195]^x[142]^x[131]^x[104]^x[76]^x[65]^x[47]^x[43]^x[42]^x[41]^x[32]^x[16]^x[15]^x[5]^x[1];
	y[14]=x[379]^x[378]^x[377]^x[376]^x[373]^x[372]^x[371]^x[370]^x[368]^x[367]^x[366]^x[365]^x[362]^x[361]^x[360]^x[359]^x[356]^x[354]^x[344]^x[335]^x[334]^x[324]^x[322]^x[282]^x[281]^x[273]^x[271]^x[262]^x[261]^x[260]^x[235]^x[224]^x[219]^x[218]^x[217]^x[216]^x[208]^x[207]^x[206]^x[205]^x[196]^x[194]^x[141]^x[130]^x[103]^x[75]^x[64]^x[46]^x[41]^x[40]^x[15]^x[14]^x[4]^x[0];
	y[13]=x[378]^x[377]^x[376]^x[375]^x[372]^x[371]^x[370]^x[369]^x[367]^x[366]^x[365]^x[364]^x[361]^x[360]^x[359]^x[358]^x[355]^x[353]^x[343]^x[334]^x[333]^x[323]^x[321]^x[281]^x[280]^x[272]^x[270]^x[261]^x[260]^x[259]^x[218]^x[217]^x[216]^x[215]^x[207]^x[206]^x[205]^x[204]^x[195]^x[193]^x[140]^x[129]^x[102]^x[45]^x[40]^x[39]^x[14]^x[13]^x[3];
	y[12]=x[377]^x[376]^x[375]^x[374]^x[371]^x[370]^x[369]^x[368]^x[366]^x[365]^x[364]^x[363]^x[360]^x[359]^x[358]^x[357]^x[354]^x[352]^x[342]^x[333]^x[332]^x[322]^x[320]^x[280]^x[279]^x[271]^x[269]^x[260]^x[259]^x[258]^x[217]^x[216]^x[215]^x[214]^x[206]^x[205]^x[204]^x[203]^x[194]^x[192]^x[101]^x[44]^x[39]^x[38]^x[13]^x[12]^x[2];
	y[11]=x[376]^x[375]^x[374]^x[370]^x[369]^x[368]^x[365]^x[363]^x[359]^x[358]^x[357]^x[352]^x[332]^x[331]^x[321]^x[279]^x[278]^x[270]^x[268]^x[259]^x[258]^x[257]^x[216]^x[215]^x[214]^x[205]^x[203]^x[192]^x[43]^x[38]^x[37]^x[12]^x[11]^x[1];
	y[10]=x[375]^x[374]^x[373]^x[369]^x[368]^x[367]^x[364]^x[363]^x[362]^x[358]^x[357]^x[356]^x[352]^x[331]^x[330]^x[320]^x[278]^x[277]^x[269]^x[267]^x[258]^x[257]^x[256]^x[215]^x[214]^x[213]^x[204]^x[203]^x[202]^x[192]^x[42]^x[37]^x[36]^x[11]^x[10]^x[0];
	y[9]=x[383]^x[382]^x[378]^x[377]^x[376]^x[374]^x[373]^x[371]^x[368]^x[367]^x[365]^x[363]^x[361]^x[357]^x[355]^x[351]^x[329]^x[287]^x[277]^x[276]^x[268]^x[257]^x[256]^x[223]^x[222]^x[214]^x[213]^x[211]^x[203]^x[201]^x[157]^x[136]^x[58]^x[41]^x[35]^x[31]^x[9];
	y[8]=x[381]^x[375]^x[373]^x[372]^x[371]^x[370]^x[367]^x[366]^x[365]^x[364]^x[362]^x[360]^x[356]^x[354]^x[350]^x[328]^x[287]^x[286]^x[276]^x[275]^x[267]^x[266]^x[256]^x[221]^x[213]^x[212]^x[211]^x[210]^x[202]^x[200]^x[156]^x[40]^x[34]^x[30]^x[8];
	y[7]=x[380]^x[374]^x[372]^x[371]^x[370]^x[369]^x[366]^x[365]^x[364]^x[363]^x[361]^x[359]^x[355]^x[353]^x[349]^x[327]^x[309]^x[298]^x[287]^x[286]^x[285]^x[275]^x[274]^x[265]^x[220]^x[212]^x[211]^x[210]^x[209]^x[201]^x[199]^x[155]^x[74]^x[68]^x[39]^x[33]^x[29]^x[7];
	y[6]=x[379]^x[373]^x[371]^x[370]^x[369]^x[368]^x[365]^x[364]^x[363]^x[362]^x[360]^x[358]^x[354]^x[352]^x[348]^x[326]^x[308]^x[297]^x[286]^x[285]^x[284]^x[274]^x[273]^x[264]^x[219]^x[211]^x[210]^x[209]^x[208]^x[200]^x[198]^x[154]^x[73]^x[67]^x[38]^x[32]^x[28]^x[6];
	y[5]=x[378]^x[374]^x[372]^x[370]^x[369]^x[367]^x[361]^x[359]^x[352]^x[347]^x[341]^x[335]^x[330]^x[325]^x[324]^x[307]^x[296]^x[285]^x[284]^x[283]^x[273]^x[272]^x[263]^x[218]^x[210]^x[209]^x[207]^x[199]^x[181]^x[170]^x[153]^x[72]^x[66]^x[54]^x[44]^x[43]^x[42]^x[37]^x[33]^x[32]^x[27]^x[5];
	y[4]=x[377]^x[371]^x[369]^x[368]^x[367]^x[366]^x[360]^x[358]^x[356]^x[346]^x[340]^x[334]^x[329]^x[324]^x[323]^x[306]^x[295]^x[284]^x[283]^x[282]^x[272]^x[271]^x[262]^x[217]^x[209]^x[208]^x[207]^x[206]^x[198]^x[196]^x[180]^x[169]^x[152]^x[71]^x[65]^x[43]^x[42]^x[41]^x[36]^x[32]^x[26]^x[4];
	y[3]=x[376]^x[370]^x[368]^x[367]^x[366]^x[365]^x[359]^x[357]^x[355]^x[345]^x[339]^x[333]^x[328]^x[323]^x[322]^x[305]^x[294]^x[283]^x[282]^x[281]^x[271]^x[270]^x[261]^x[216]^x[208]^x[207]^x[206]^x[205]^x[197]^x[195]^x[179]^x[168]^x[151]^x[70]^x[64]^x[42]^x[41]^x[40]^x[35]^x[25]^x[3];
	y[2]=x[375]^x[369]^x[367]^x[366]^x[365]^x[364]^x[358]^x[356]^x[354]^x[344]^x[338]^x[332]^x[327]^x[322]^x[321]^x[304]^x[293]^x[282]^x[281]^x[280]^x[270]^x[269]^x[260]^x[215]^x[207]^x[206]^x[205]^x[204]^x[196]^x[194]^x[178]^x[167]^x[150]^x[69]^x[41]^x[40]^x[39]^x[34]^x[24]^x[2];
	y[1]=x[374]^x[368]^x[366]^x[365]^x[364]^x[363]^x[357]^x[355]^x[353]^x[343]^x[337]^x[331]^x[326]^x[321]^x[320]^x[281]^x[280]^x[279]^x[269]^x[268]^x[259]^x[214]^x[206]^x[205]^x[204]^x[203]^x[195]^x[193]^x[177]^x[166]^x[40]^x[39]^x[38]^x[33]^x[23]^x[1];
	y[0]=x[374]^x[368]^x[365]^x[364]^x[363]^x[357]^x[354]^x[342]^x[336]^x[325]^x[320]^x[280]^x[279]^x[278]^x[268]^x[267]^x[258]^x[214]^x[205]^x[204]^x[203]^x[194]^x[176]^x[165]^x[39]^x[38]^x[37]^x[32]^x[22]^x[0];
	return y;
endfunction

(* noinline *)
function Bit#(384) update_state(Bit#(384) x);
	Bit#(384) x_new = 0;
	x_new[383]=x[383]^x[373]^x[363]^x[352]^x[346]^x[345]^x[336]^x[334]^x[325]^x[319]^x[318]^x[309]^x[307]^x[298]^x[285]^x[282]^x[279]^x[278]^x[276]^x[274]^x[272]^x[270]^x[268]^x[267]^x[266]^x[263]^x[261]^x[260]^x[257]^x[255]^x[247]^x[246]^x[245]^x[235]^x[234]^x[225]^x[191]^x[186]^x[181]^x[176]^x[170]^x[165]^x[125]^x[122]^x[118]^x[114]^x[110]^x[107]^x[106]^x[104]^x[103]^x[95]^x[89]^x[83]^x[77]^x[49]^x[31]^x[26]^x[25]^x[16]^x[12]^x[11]^x[6]^x[1];
	x_new[382]=x[383]^x[382]^x[372]^x[318]^x[317]^x[308]^x[306]^x[297]^x[286]^x[284]^x[280]^x[278]^x[277]^x[274]^x[273]^x[271]^x[268]^x[267]^x[266]^x[265]^x[263]^x[262]^x[260]^x[259]^x[257]^x[256]^x[254]^x[246]^x[245]^x[244]^x[234]^x[233]^x[224]^x[126]^x[124]^x[117]^x[114]^x[113]^x[106]^x[105]^x[103]^x[102]^x[94]^x[88]^x[82]^x[76]^x[48]^x[30]^x[24]^x[11]^x[10]^x[5]^x[4]^x[0];
	x_new[381]=x[382]^x[381]^x[371]^x[317]^x[316]^x[307]^x[305]^x[296]^x[285]^x[283]^x[279]^x[277]^x[276]^x[273]^x[272]^x[270]^x[266]^x[265]^x[264]^x[262]^x[261]^x[259]^x[258]^x[255]^x[253]^x[245]^x[244]^x[243]^x[234]^x[233]^x[232]^x[125]^x[123]^x[116]^x[113]^x[112]^x[105]^x[104]^x[102]^x[101]^x[93]^x[87]^x[81]^x[75]^x[47]^x[31]^x[29]^x[25]^x[23]^x[9]^x[3];
	x_new[380]=x[381]^x[380]^x[370]^x[316]^x[315]^x[306]^x[304]^x[295]^x[284]^x[282]^x[278]^x[276]^x[275]^x[272]^x[271]^x[269]^x[265]^x[264]^x[263]^x[261]^x[260]^x[258]^x[257]^x[254]^x[252]^x[244]^x[243]^x[242]^x[233]^x[232]^x[231]^x[124]^x[122]^x[115]^x[112]^x[111]^x[104]^x[103]^x[101]^x[100]^x[92]^x[86]^x[80]^x[74]^x[46]^x[30]^x[28]^x[24]^x[22]^x[8]^x[2];
	x_new[379]=x[380]^x[379]^x[369]^x[315]^x[314]^x[305]^x[303]^x[294]^x[283]^x[281]^x[277]^x[275]^x[274]^x[271]^x[270]^x[268]^x[264]^x[263]^x[262]^x[260]^x[259]^x[257]^x[256]^x[253]^x[251]^x[243]^x[242]^x[241]^x[232]^x[231]^x[230]^x[123]^x[121]^x[114]^x[111]^x[110]^x[103]^x[102]^x[100]^x[99]^x[91]^x[85]^x[79]^x[73]^x[45]^x[29]^x[27]^x[23]^x[21]^x[7]^x[1];
	x_new[378]=x[379]^x[378]^x[368]^x[351]^x[350]^x[341]^x[340]^x[339]^x[331]^x[320]^x[314]^x[313]^x[304]^x[302]^x[293]^x[285]^x[282]^x[280]^x[277]^x[275]^x[274]^x[273]^x[270]^x[269]^x[267]^x[265]^x[262]^x[261]^x[259]^x[258]^x[256]^x[252]^x[250]^x[242]^x[241]^x[240]^x[231]^x[230]^x[229]^x[186]^x[181]^x[175]^x[171]^x[160]^x[159]^x[138]^x[122]^x[120]^x[117]^x[116]^x[115]^x[113]^x[111]^x[102]^x[101]^x[99]^x[98]^x[90]^x[84]^x[78]^x[72]^x[44]^x[28]^x[26]^x[22]^x[21]^x[20]^x[11]^x[6];
	x_new[377]=x[378]^x[377]^x[367]^x[349]^x[340]^x[338]^x[313]^x[312]^x[303]^x[301]^x[292]^x[287]^x[284]^x[281]^x[279]^x[276]^x[274]^x[273]^x[272]^x[269]^x[268]^x[264]^x[261]^x[260]^x[258]^x[257]^x[251]^x[249]^x[241]^x[240]^x[239]^x[230]^x[229]^x[228]^x[180]^x[174]^x[158]^x[137]^x[127]^x[119]^x[116]^x[114]^x[112]^x[110]^x[109]^x[106]^x[101]^x[98]^x[97]^x[89]^x[83]^x[77]^x[71]^x[43]^x[27]^x[25]^x[21]^x[20]^x[19]^x[5];
	x_new[376]=x[377]^x[376]^x[366]^x[348]^x[339]^x[337]^x[312]^x[311]^x[302]^x[300]^x[291]^x[286]^x[283]^x[280]^x[278]^x[275]^x[273]^x[272]^x[271]^x[268]^x[267]^x[263]^x[260]^x[259]^x[257]^x[256]^x[250]^x[248]^x[240]^x[239]^x[238]^x[229]^x[228]^x[227]^x[179]^x[173]^x[157]^x[136]^x[126]^x[118]^x[115]^x[113]^x[111]^x[109]^x[108]^x[105]^x[100]^x[97]^x[96]^x[88]^x[82]^x[76]^x[70]^x[42]^x[26]^x[24]^x[20]^x[19]^x[18]^x[4];
	x_new[375]=x[376]^x[375]^x[365]^x[347]^x[338]^x[336]^x[311]^x[310]^x[301]^x[299]^x[290]^x[285]^x[282]^x[279]^x[274]^x[272]^x[270]^x[262]^x[260]^x[259]^x[258]^x[249]^x[247]^x[239]^x[238]^x[237]^x[228]^x[227]^x[226]^x[178]^x[172]^x[156]^x[135]^x[125]^x[114]^x[112]^x[110]^x[108]^x[106]^x[104]^x[99]^x[87]^x[81]^x[75]^x[69]^x[41]^x[25]^x[23]^x[19]^x[18]^x[17]^x[3];
	x_new[374]=x[375]^x[374]^x[364]^x[346]^x[337]^x[335]^x[310]^x[309]^x[300]^x[298]^x[289]^x[284]^x[281]^x[278]^x[273]^x[271]^x[269]^x[261]^x[259]^x[258]^x[257]^x[248]^x[246]^x[238]^x[237]^x[236]^x[227]^x[226]^x[225]^x[177]^x[171]^x[155]^x[134]^x[124]^x[113]^x[111]^x[109]^x[107]^x[105]^x[103]^x[98]^x[86]^x[80]^x[74]^x[68]^x[40]^x[24]^x[22]^x[18]^x[17]^x[16]^x[2];
	x_new[373]=x[374]^x[373]^x[363]^x[345]^x[336]^x[334]^x[309]^x[308]^x[299]^x[297]^x[288]^x[283]^x[280]^x[272]^x[271]^x[270]^x[268]^x[266]^x[258]^x[257]^x[256]^x[247]^x[245]^x[237]^x[236]^x[235]^x[226]^x[225]^x[224]^x[176]^x[171]^x[160]^x[154]^x[133]^x[123]^x[117]^x[112]^x[110]^x[108]^x[104]^x[102]^x[97]^x[85]^x[79]^x[73]^x[67]^x[39]^x[23]^x[21]^x[17]^x[16]^x[15]^x[1];
	x_new[372]=x[373]^x[372]^x[362]^x[346]^x[345]^x[334]^x[319]^x[308]^x[307]^x[296]^x[287]^x[286]^x[285]^x[282]^x[281]^x[280]^x[279]^x[276]^x[274]^x[270]^x[268]^x[267]^x[266]^x[260]^x[256]^x[255]^x[246]^x[244]^x[236]^x[235]^x[225]^x[224]^x[191]^x[190]^x[186]^x[169]^x[127]^x[126]^x[125]^x[122]^x[114]^x[110]^x[107]^x[106]^x[104]^x[101]^x[96]^x[84]^x[78]^x[72]^x[66]^x[38]^x[26]^x[22]^x[20]^x[16]^x[14]^x[0];
	x_new[371]=x[372]^x[371]^x[361]^x[318]^x[307]^x[306]^x[295]^x[287]^x[286]^x[285]^x[284]^x[281]^x[280]^x[279]^x[278]^x[275]^x[273]^x[269]^x[267]^x[265]^x[259]^x[255]^x[254]^x[245]^x[243]^x[235]^x[224]^x[189]^x[179]^x[168]^x[127]^x[126]^x[125]^x[124]^x[115]^x[113]^x[105]^x[83]^x[77]^x[71]^x[65]^x[37]^x[31]^x[25]^x[21]^x[19]^x[15]^x[13]^x[10]^x[4];
	x_new[370]=x[371]^x[370]^x[360]^x[317]^x[306]^x[305]^x[294]^x[286]^x[285]^x[284]^x[283]^x[280]^x[279]^x[278]^x[277]^x[274]^x[272]^x[268]^x[266]^x[264]^x[258]^x[255]^x[254]^x[253]^x[244]^x[242]^x[188]^x[178]^x[167]^x[126]^x[125]^x[124]^x[123]^x[114]^x[112]^x[104]^x[82]^x[76]^x[70]^x[64]^x[36]^x[30]^x[24]^x[20]^x[18]^x[14]^x[12]^x[9]^x[3];
	x_new[369]=x[370]^x[369]^x[359]^x[342]^x[341]^x[330]^x[320]^x[316]^x[305]^x[304]^x[293]^x[285]^x[284]^x[283]^x[282]^x[279]^x[278]^x[277]^x[276]^x[273]^x[271]^x[266]^x[265]^x[263]^x[257]^x[256]^x[254]^x[253]^x[252]^x[243]^x[241]^x[187]^x[177]^x[166]^x[125]^x[124]^x[123]^x[122]^x[113]^x[111]^x[107]^x[106]^x[103]^x[101]^x[100]^x[96]^x[81]^x[75]^x[69]^x[35]^x[29]^x[23]^x[19]^x[17]^x[13]^x[11]^x[8]^x[2];
	x_new[368]=x[369]^x[368]^x[358]^x[340]^x[329]^x[315]^x[304]^x[303]^x[292]^x[284]^x[283]^x[282]^x[281]^x[278]^x[277]^x[276]^x[275]^x[272]^x[270]^x[266]^x[265]^x[264]^x[262]^x[256]^x[253]^x[252]^x[251]^x[242]^x[240]^x[186]^x[176]^x[165]^x[124]^x[123]^x[122]^x[121]^x[112]^x[110]^x[105]^x[102]^x[99]^x[80]^x[74]^x[68]^x[34]^x[28]^x[22]^x[18]^x[16]^x[12]^x[10]^x[7]^x[1];
	x_new[367]=x[368]^x[367]^x[357]^x[341]^x[339]^x[330]^x[328]^x[314]^x[303]^x[302]^x[291]^x[283]^x[282]^x[281]^x[280]^x[277]^x[276]^x[275]^x[274]^x[271]^x[269]^x[266]^x[265]^x[264]^x[263]^x[261]^x[252]^x[251]^x[250]^x[241]^x[239]^x[185]^x[181]^x[170]^x[123]^x[122]^x[121]^x[120]^x[111]^x[109]^x[106]^x[104]^x[101]^x[100]^x[98]^x[79]^x[73]^x[67]^x[33]^x[27]^x[17]^x[15]^x[11]^x[10]^x[9]^x[6]^x[0];
	x_new[366]=x[367]^x[366]^x[356]^x[340]^x[338]^x[329]^x[327]^x[313]^x[302]^x[301]^x[290]^x[282]^x[281]^x[280]^x[279]^x[276]^x[275]^x[274]^x[273]^x[270]^x[268]^x[265]^x[264]^x[263]^x[262]^x[260]^x[251]^x[250]^x[249]^x[240]^x[238]^x[184]^x[180]^x[169]^x[122]^x[121]^x[120]^x[119]^x[110]^x[108]^x[105]^x[103]^x[100]^x[99]^x[97]^x[78]^x[72]^x[66]^x[32]^x[26]^x[16]^x[14]^x[10]^x[9]^x[8]^x[5];
	x_new[365]=x[366]^x[365]^x[355]^x[339]^x[337]^x[328]^x[326]^x[312]^x[301]^x[300]^x[289]^x[281]^x[280]^x[279]^x[278]^x[275]^x[274]^x[273]^x[272]^x[269]^x[267]^x[264]^x[263]^x[262]^x[261]^x[259]^x[250]^x[249]^x[248]^x[239]^x[237]^x[183]^x[179]^x[168]^x[121]^x[120]^x[119]^x[118]^x[109]^x[107]^x[104]^x[102]^x[99]^x[98]^x[96]^x[77]^x[71]^x[65]^x[25]^x[15]^x[13]^x[9]^x[8]^x[7]^x[4];
	x_new[364]=x[365]^x[364]^x[354]^x[338]^x[336]^x[327]^x[325]^x[311]^x[300]^x[299]^x[288]^x[280]^x[279]^x[278]^x[274]^x[273]^x[272]^x[268]^x[263]^x[262]^x[261]^x[258]^x[249]^x[248]^x[247]^x[238]^x[236]^x[182]^x[178]^x[167]^x[120]^x[119]^x[118]^x[108]^x[103]^x[101]^x[98]^x[97]^x[76]^x[70]^x[64]^x[24]^x[14]^x[12]^x[8]^x[7]^x[6]^x[3];
	x_new[363]=x[364]^x[363]^x[353]^x[337]^x[336]^x[326]^x[325]^x[310]^x[299]^x[279]^x[278]^x[273]^x[272]^x[262]^x[261]^x[257]^x[256]^x[248]^x[247]^x[246]^x[237]^x[235]^x[182]^x[177]^x[171]^x[166]^x[119]^x[118]^x[102]^x[101]^x[97]^x[75]^x[69]^x[23]^x[13]^x[11]^x[7]^x[6]^x[5]^x[2];
	x_new[362]=x[363]^x[362]^x[352]^x[336]^x[325]^x[309]^x[298]^x[278]^x[277]^x[272]^x[271]^x[266]^x[261]^x[260]^x[256]^x[247]^x[246]^x[245]^x[236]^x[234]^x[176]^x[165]^x[118]^x[117]^x[106]^x[101]^x[96]^x[74]^x[68]^x[22]^x[12]^x[10]^x[6]^x[5]^x[4]^x[1];
	x_new[361]=x[383]^x[361]^x[308]^x[297]^x[287]^x[286]^x[281]^x[280]^x[277]^x[276]^x[275]^x[274]^x[271]^x[270]^x[269]^x[268]^x[266]^x[265]^x[263]^x[260]^x[259]^x[257]^x[246]^x[245]^x[244]^x[235]^x[233]^x[180]^x[179]^x[169]^x[127]^x[126]^x[117]^x[116]^x[115]^x[114]^x[106]^x[105]^x[103]^x[73]^x[67]^x[21]^x[15]^x[11]^x[9]^x[5]^x[3]^x[0];
	x_new[360]=x[382]^x[360]^x[307]^x[296]^x[286]^x[285]^x[280]^x[279]^x[276]^x[275]^x[274]^x[273]^x[270]^x[269]^x[268]^x[267]^x[265]^x[264]^x[262]^x[259]^x[258]^x[256]^x[245]^x[244]^x[243]^x[234]^x[232]^x[179]^x[178]^x[168]^x[126]^x[125]^x[116]^x[115]^x[114]^x[113]^x[105]^x[104]^x[102]^x[72]^x[66]^x[31]^x[25]^x[20]^x[14]^x[8]^x[2];
	x_new[359]=x[381]^x[359]^x[306]^x[295]^x[285]^x[284]^x[279]^x[278]^x[275]^x[274]^x[273]^x[272]^x[269]^x[268]^x[267]^x[264]^x[263]^x[261]^x[258]^x[257]^x[244]^x[243]^x[242]^x[233]^x[231]^x[178]^x[177]^x[167]^x[125]^x[124]^x[115]^x[114]^x[113]^x[112]^x[104]^x[103]^x[101]^x[71]^x[65]^x[30]^x[24]^x[19]^x[13]^x[7]^x[1];
	x_new[358]=x[380]^x[358]^x[305]^x[294]^x[284]^x[283]^x[278]^x[277]^x[274]^x[273]^x[272]^x[271]^x[268]^x[267]^x[266]^x[263]^x[262]^x[260]^x[257]^x[256]^x[243]^x[242]^x[241]^x[232]^x[230]^x[177]^x[176]^x[166]^x[124]^x[123]^x[114]^x[113]^x[112]^x[111]^x[103]^x[102]^x[100]^x[70]^x[64]^x[29]^x[23]^x[18]^x[12]^x[6]^x[0];
	x_new[357]=x[379]^x[357]^x[342]^x[320]^x[304]^x[293]^x[283]^x[282]^x[277]^x[276]^x[273]^x[272]^x[271]^x[270]^x[266]^x[265]^x[262]^x[261]^x[259]^x[242]^x[241]^x[240]^x[231]^x[229]^x[182]^x[175]^x[160]^x[138]^x[123]^x[122]^x[113]^x[112]^x[111]^x[110]^x[107]^x[102]^x[99]^x[96]^x[69]^x[28]^x[17]^x[11]^x[5]^x[0];
	x_new[356]=x[378]^x[356]^x[341]^x[330]^x[303]^x[292]^x[282]^x[281]^x[276]^x[275]^x[272]^x[271]^x[270]^x[269]^x[265]^x[264]^x[261]^x[260]^x[258]^x[241]^x[240]^x[239]^x[230]^x[228]^x[181]^x[174]^x[170]^x[137]^x[122]^x[121]^x[112]^x[111]^x[110]^x[109]^x[106]^x[101]^x[98]^x[68]^x[27]^x[16]^x[4];
	x_new[355]=x[377]^x[355]^x[340]^x[329]^x[302]^x[291]^x[281]^x[280]^x[275]^x[274]^x[271]^x[270]^x[269]^x[268]^x[264]^x[263]^x[260]^x[259]^x[257]^x[240]^x[239]^x[238]^x[229]^x[227]^x[180]^x[173]^x[169]^x[136]^x[121]^x[120]^x[111]^x[110]^x[109]^x[108]^x[105]^x[100]^x[97]^x[67]^x[26]^x[15]^x[3];
	x_new[354]=x[376]^x[354]^x[339]^x[328]^x[301]^x[290]^x[280]^x[279]^x[274]^x[273]^x[270]^x[269]^x[268]^x[267]^x[263]^x[262]^x[259]^x[258]^x[256]^x[239]^x[238]^x[237]^x[228]^x[226]^x[179]^x[172]^x[168]^x[135]^x[120]^x[119]^x[110]^x[109]^x[108]^x[107]^x[104]^x[99]^x[96]^x[66]^x[25]^x[14]^x[2];
	x_new[353]=x[375]^x[353]^x[338]^x[327]^x[300]^x[289]^x[279]^x[278]^x[273]^x[272]^x[269]^x[268]^x[267]^x[262]^x[261]^x[258]^x[257]^x[238]^x[237]^x[236]^x[227]^x[225]^x[178]^x[171]^x[167]^x[134]^x[119]^x[118]^x[109]^x[108]^x[107]^x[103]^x[98]^x[65]^x[24]^x[13]^x[1];
	x_new[352]=x[374]^x[352]^x[337]^x[326]^x[299]^x[288]^x[278]^x[272]^x[268]^x[267]^x[261]^x[257]^x[256]^x[237]^x[236]^x[235]^x[226]^x[224]^x[177]^x[171]^x[166]^x[160]^x[133]^x[118]^x[108]^x[107]^x[102]^x[97]^x[64]^x[23]^x[12]^x[0];
	x_new[351]=x[383]^x[379]^x[378]^x[377]^x[375]^x[374]^x[373]^x[369]^x[367]^x[363]^x[362]^x[358]^x[357]^x[356]^x[353]^x[351]^x[341]^x[331]^x[320]^x[314]^x[313]^x[304]^x[302]^x[293]^x[287]^x[286]^x[277]^x[275]^x[266]^x[253]^x[250]^x[247]^x[246]^x[244]^x[242]^x[240]^x[238]^x[236]^x[235]^x[234]^x[231]^x[229]^x[228]^x[225]^x[223]^x[215]^x[214]^x[213]^x[203]^x[202]^x[193]^x[149]^x[148]^x[147]^x[140]^x[139]^x[129]^x[128]^x[93]^x[90]^x[86]^x[82]^x[78]^x[75]^x[74]^x[72]^x[71]^x[63]^x[57]^x[51]^x[45]^x[17];
	x_new[350]=x[382]^x[376]^x[374]^x[373]^x[372]^x[368]^x[367]^x[366]^x[362]^x[361]^x[357]^x[356]^x[355]^x[352]^x[351]^x[350]^x[340]^x[286]^x[285]^x[276]^x[274]^x[265]^x[254]^x[252]^x[248]^x[246]^x[245]^x[242]^x[241]^x[239]^x[236]^x[235]^x[234]^x[233]^x[231]^x[230]^x[228]^x[227]^x[225]^x[224]^x[222]^x[214]^x[213]^x[212]^x[202]^x[201]^x[192]^x[158]^x[146]^x[139]^x[138]^x[128]^x[94]^x[92]^x[85]^x[82]^x[81]^x[74]^x[73]^x[71]^x[70]^x[62]^x[56]^x[50]^x[44]^x[16];
	x_new[349]=x[383]^x[381]^x[377]^x[375]^x[373]^x[372]^x[371]^x[367]^x[366]^x[365]^x[362]^x[361]^x[360]^x[356]^x[355]^x[354]^x[350]^x[349]^x[339]^x[285]^x[284]^x[275]^x[273]^x[264]^x[253]^x[251]^x[247]^x[245]^x[244]^x[241]^x[240]^x[238]^x[234]^x[233]^x[232]^x[230]^x[229]^x[227]^x[226]^x[223]^x[221]^x[213]^x[212]^x[211]^x[202]^x[201]^x[200]^x[159]^x[157]^x[147]^x[145]^x[137]^x[93]^x[91]^x[84]^x[81]^x[80]^x[73]^x[72]^x[70]^x[69]^x[61]^x[55]^x[49]^x[43]^x[15];
	x_new[348]=x[382]^x[380]^x[376]^x[374]^x[372]^x[371]^x[370]^x[366]^x[365]^x[364]^x[361]^x[360]^x[359]^x[355]^x[354]^x[353]^x[349]^x[348]^x[338]^x[284]^x[283]^x[274]^x[272]^x[263]^x[252]^x[250]^x[246]^x[244]^x[243]^x[240]^x[239]^x[237]^x[233]^x[232]^x[231]^x[229]^x[228]^x[226]^x[225]^x[222]^x[220]^x[212]^x[211]^x[210]^x[201]^x[200]^x[199]^x[158]^x[156]^x[146]^x[144]^x[136]^x[92]^x[90]^x[83]^x[80]^x[79]^x[72]^x[71]^x[69]^x[68]^x[60]^x[54]^x[48]^x[42]^x[14];
	x_new[347]=x[381]^x[379]^x[375]^x[373]^x[371]^x[370]^x[369]^x[365]^x[364]^x[363]^x[360]^x[359]^x[358]^x[354]^x[353]^x[352]^x[348]^x[347]^x[337]^x[283]^x[282]^x[273]^x[271]^x[262]^x[251]^x[249]^x[245]^x[243]^x[242]^x[239]^x[238]^x[236]^x[232]^x[231]^x[230]^x[228]^x[227]^x[225]^x[224]^x[221]^x[219]^x[211]^x[210]^x[209]^x[200]^x[199]^x[198]^x[157]^x[155]^x[145]^x[143]^x[135]^x[91]^x[89]^x[82]^x[79]^x[78]^x[71]^x[70]^x[68]^x[67]^x[59]^x[53]^x[47]^x[41]^x[13];
	x_new[346]=x[383]^x[380]^x[378]^x[373]^x[372]^x[370]^x[369]^x[368]^x[364]^x[359]^x[358]^x[357]^x[353]^x[352]^x[347]^x[346]^x[336]^x[319]^x[318]^x[309]^x[308]^x[307]^x[299]^x[288]^x[282]^x[281]^x[272]^x[270]^x[261]^x[253]^x[250]^x[248]^x[245]^x[243]^x[242]^x[241]^x[238]^x[237]^x[235]^x[233]^x[230]^x[229]^x[227]^x[226]^x[224]^x[220]^x[218]^x[210]^x[209]^x[208]^x[199]^x[198]^x[197]^x[156]^x[144]^x[142]^x[134]^x[133]^x[127]^x[106]^x[90]^x[88]^x[85]^x[84]^x[83]^x[81]^x[79]^x[70]^x[69]^x[67]^x[66]^x[58]^x[52]^x[46]^x[40]^x[12];
	x_new[345]=x[383]^x[382]^x[379]^x[377]^x[373]^x[372]^x[371]^x[369]^x[368]^x[367]^x[363]^x[358]^x[357]^x[356]^x[352]^x[346]^x[345]^x[335]^x[317]^x[308]^x[306]^x[281]^x[280]^x[271]^x[269]^x[260]^x[255]^x[252]^x[249]^x[247]^x[244]^x[242]^x[241]^x[240]^x[237]^x[236]^x[232]^x[229]^x[228]^x[226]^x[225]^x[219]^x[217]^x[209]^x[208]^x[207]^x[198]^x[197]^x[196]^x[155]^x[153]^x[143]^x[141]^x[133]^x[126]^x[105]^x[95]^x[87]^x[84]^x[82]^x[80]^x[78]^x[77]^x[74]^x[69]^x[66]^x[65]^x[57]^x[51]^x[45]^x[39]^x[11];
	x_new[344]=x[383]^x[382]^x[381]^x[378]^x[376]^x[372]^x[371]^x[370]^x[368]^x[367]^x[366]^x[357]^x[356]^x[355]^x[345]^x[344]^x[334]^x[316]^x[307]^x[305]^x[280]^x[279]^x[270]^x[268]^x[259]^x[254]^x[251]^x[248]^x[246]^x[243]^x[241]^x[240]^x[239]^x[236]^x[235]^x[231]^x[228]^x[227]^x[225]^x[224]^x[218]^x[216]^x[208]^x[207]^x[206]^x[197]^x[196]^x[195]^x[154]^x[152]^x[142]^x[140]^x[132]^x[125]^x[104]^x[94]^x[86]^x[83]^x[81]^x[79]^x[77]^x[76]^x[73]^x[68]^x[65]^x[64]^x[56]^x[50]^x[44]^x[38]^x[10];
	x_new[343]=x[382]^x[381]^x[380]^x[377]^x[375]^x[371]^x[370]^x[369]^x[367]^x[366]^x[365]^x[356]^x[355]^x[354]^x[344]^x[343]^x[333]^x[315]^x[306]^x[304]^x[279]^x[278]^x[269]^x[267]^x[258]^x[253]^x[250]^x[247]^x[242]^x[240]^x[238]^x[230]^x[228]^x[227]^x[226]^x[217]^x[215]^x[207]^x[206]^x[205]^x[196]^x[195]^x[194]^x[153]^x[151]^x[141]^x[139]^x[131]^x[124]^x[103]^x[93]^x[82]^x[80]^x[78]^x[76]^x[74]^x[72]^x[67]^x[55]^x[49]^x[43]^x[37]^x[9];
	x_new[342]=x[381]^x[380]^x[379]^x[376]^x[374]^x[370]^x[369]^x[368]^x[366]^x[365]^x[364]^x[355]^x[354]^x[353]^x[343]^x[342]^x[332]^x[314]^x[305]^x[303]^x[278]^x[277]^x[268]^x[266]^x[257]^x[252]^x[249]^x[246]^x[241]^x[239]^x[237]^x[229]^x[227]^x[226]^x[225]^x[216]^x[214]^x[206]^x[205]^x[204]^x[195]^x[194]^x[193]^x[152]^x[150]^x[140]^x[138]^x[130]^x[123]^x[102]^x[92]^x[81]^x[79]^x[77]^x[75]^x[73]^x[71]^x[66]^x[54]^x[48]^x[42]^x[36]^x[8];
	x_new[341]=x[380]^x[379]^x[378]^x[375]^x[373]^x[369]^x[368]^x[367]^x[365]^x[364]^x[363]^x[354]^x[353]^x[352]^x[342]^x[341]^x[331]^x[313]^x[304]^x[302]^x[277]^x[276]^x[267]^x[265]^x[256]^x[251]^x[248]^x[240]^x[239]^x[238]^x[236]^x[234]^x[226]^x[225]^x[224]^x[215]^x[213]^x[205]^x[204]^x[203]^x[194]^x[193]^x[192]^x[151]^x[149]^x[138]^x[137]^x[129]^x[128]^x[122]^x[101]^x[91]^x[85]^x[80]^x[78]^x[76]^x[72]^x[70]^x[65]^x[53]^x[47]^x[41]^x[35]^x[7];
	x_new[340]=x[383]^x[379]^x[378]^x[377]^x[374]^x[372]^x[366]^x[364]^x[363]^x[357]^x[353]^x[352]^x[341]^x[340]^x[330]^x[314]^x[313]^x[302]^x[287]^x[276]^x[275]^x[264]^x[255]^x[254]^x[253]^x[250]^x[249]^x[248]^x[247]^x[244]^x[242]^x[238]^x[236]^x[235]^x[234]^x[228]^x[224]^x[223]^x[214]^x[212]^x[204]^x[203]^x[193]^x[192]^x[159]^x[158]^x[150]^x[138]^x[137]^x[136]^x[128]^x[95]^x[94]^x[93]^x[90]^x[82]^x[78]^x[75]^x[74]^x[72]^x[69]^x[64]^x[52]^x[46]^x[40]^x[34]^x[6];
	x_new[339]=x[383]^x[382]^x[378]^x[377]^x[376]^x[373]^x[371]^x[367]^x[365]^x[363]^x[352]^x[340]^x[339]^x[329]^x[286]^x[275]^x[274]^x[263]^x[255]^x[254]^x[253]^x[252]^x[249]^x[248]^x[247]^x[246]^x[243]^x[241]^x[237]^x[235]^x[233]^x[227]^x[223]^x[222]^x[213]^x[211]^x[203]^x[192]^x[159]^x[157]^x[149]^x[147]^x[138]^x[137]^x[136]^x[135]^x[95]^x[94]^x[93]^x[92]^x[83]^x[81]^x[73]^x[51]^x[45]^x[39]^x[33]^x[5];
	x_new[338]=x[383]^x[382]^x[381]^x[377]^x[376]^x[375]^x[372]^x[370]^x[366]^x[364]^x[339]^x[338]^x[328]^x[285]^x[274]^x[273]^x[262]^x[254]^x[253]^x[252]^x[251]^x[248]^x[247]^x[246]^x[245]^x[242]^x[240]^x[236]^x[234]^x[232]^x[226]^x[223]^x[222]^x[221]^x[212]^x[210]^x[158]^x[156]^x[148]^x[146]^x[137]^x[136]^x[135]^x[134]^x[94]^x[93]^x[92]^x[91]^x[82]^x[80]^x[72]^x[50]^x[44]^x[38]^x[32]^x[4];
	x_new[337]=x[382]^x[381]^x[380]^x[376]^x[375]^x[374]^x[371]^x[369]^x[365]^x[363]^x[338]^x[337]^x[327]^x[310]^x[309]^x[298]^x[288]^x[284]^x[273]^x[272]^x[261]^x[253]^x[252]^x[251]^x[250]^x[247]^x[246]^x[245]^x[244]^x[241]^x[239]^x[234]^x[233]^x[231]^x[225]^x[224]^x[222]^x[221]^x[220]^x[211]^x[209]^x[157]^x[155]^x[147]^x[145]^x[136]^x[135]^x[134]^x[133]^x[93]^x[92]^x[91]^x[90]^x[81]^x[79]^x[75]^x[74]^x[71]^x[69]^x[68]^x[64]^x[49]^x[43]^x[37]^x[3];
	x_new[336]=x[381]^x[380]^x[379]^x[375]^x[374]^x[373]^x[370]^x[368]^x[364]^x[362]^x[337]^x[336]^x[326]^x[308]^x[297]^x[283]^x[272]^x[271]^x[260]^x[252]^x[251]^x[250]^x[249]^x[246]^x[245]^x[244]^x[243]^x[240]^x[238]^x[234]^x[233]^x[232]^x[230]^x[224]^x[221]^x[220]^x[219]^x[210]^x[208]^x[156]^x[154]^x[146]^x[144]^x[135]^x[134]^x[133]^x[132]^x[92]^x[91]^x[90]^x[89]^x[80]^x[78]^x[73]^x[70]^x[67]^x[48]^x[42]^x[36]^x[2];
	x_new[335]=x[380]^x[379]^x[378]^x[374]^x[373]^x[372]^x[369]^x[367]^x[362]^x[361]^x[352]^x[336]^x[335]^x[325]^x[309]^x[307]^x[298]^x[296]^x[282]^x[271]^x[270]^x[259]^x[251]^x[250]^x[249]^x[248]^x[245]^x[244]^x[243]^x[242]^x[239]^x[237]^x[234]^x[233]^x[232]^x[231]^x[229]^x[220]^x[219]^x[218]^x[209]^x[207]^x[155]^x[153]^x[145]^x[143]^x[134]^x[133]^x[132]^x[131]^x[91]^x[90]^x[89]^x[88]^x[79]^x[77]^x[74]^x[72]^x[69]^x[68]^x[66]^x[47]^x[41]^x[35]^x[1];
	x_new[334]=x[379]^x[378]^x[377]^x[373]^x[372]^x[371]^x[368]^x[366]^x[362]^x[361]^x[360]^x[335]^x[334]^x[324]^x[308]^x[306]^x[297]^x[295]^x[281]^x[270]^x[269]^x[258]^x[250]^x[249]^x[248]^x[247]^x[244]^x[243]^x[242]^x[241]^x[238]^x[236]^x[233]^x[232]^x[231]^x[230]^x[228]^x[219]^x[218]^x[217]^x[208]^x[206]^x[154]^x[152]^x[144]^x[142]^x[133]^x[132]^x[131]^x[130]^x[90]^x[89]^x[88]^x[87]^x[78]^x[76]^x[73]^x[71]^x[68]^x[67]^x[65]^x[46]^x[40]^x[34]^x[0];
	x_new[333]=x[378]^x[377]^x[376]^x[372]^x[371]^x[370]^x[367]^x[365]^x[361]^x[360]^x[359]^x[334]^x[333]^x[323]^x[307]^x[305]^x[296]^x[294]^x[280]^x[269]^x[268]^x[257]^x[249]^x[248]^x[247]^x[246]^x[243]^x[242]^x[241]^x[240]^x[237]^x[235]^x[232]^x[231]^x[230]^x[229]^x[227]^x[218]^x[217]^x[216]^x[207]^x[205]^x[153]^x[151]^x[143]^x[141]^x[132]^x[131]^x[130]^x[129]^x[89]^x[88]^x[87]^x[86]^x[77]^x[75]^x[72]^x[70]^x[67]^x[66]^x[64]^x[45]^x[39]^x[33];
	x_new[332]=x[377]^x[376]^x[375]^x[371]^x[370]^x[369]^x[366]^x[364]^x[360]^x[359]^x[358]^x[333]^x[332]^x[322]^x[306]^x[304]^x[295]^x[293]^x[279]^x[268]^x[267]^x[256]^x[248]^x[247]^x[246]^x[242]^x[241]^x[240]^x[236]^x[231]^x[230]^x[229]^x[226]^x[217]^x[216]^x[215]^x[206]^x[204]^x[152]^x[150]^x[142]^x[140]^x[131]^x[130]^x[129]^x[128]^x[88]^x[87]^x[86]^x[76]^x[71]^x[69]^x[66]^x[65]^x[44]^x[38]^x[32];
	x_new[331]=x[376]^x[375]^x[374]^x[370]^x[369]^x[368]^x[365]^x[363]^x[359]^x[358]^x[357]^x[332]^x[331]^x[321]^x[305]^x[304]^x[294]^x[293]^x[278]^x[267]^x[247]^x[246]^x[241]^x[240]^x[230]^x[229]^x[225]^x[224]^x[216]^x[215]^x[214]^x[205]^x[203]^x[151]^x[150]^x[141]^x[130]^x[129]^x[128]^x[87]^x[86]^x[70]^x[69]^x[65]^x[43]^x[37];
	x_new[330]=x[375]^x[374]^x[373]^x[369]^x[368]^x[367]^x[364]^x[362]^x[358]^x[357]^x[356]^x[331]^x[330]^x[320]^x[304]^x[293]^x[277]^x[266]^x[246]^x[245]^x[240]^x[239]^x[234]^x[229]^x[228]^x[224]^x[215]^x[214]^x[213]^x[204]^x[202]^x[150]^x[140]^x[138]^x[129]^x[128]^x[86]^x[85]^x[74]^x[69]^x[64]^x[42]^x[36];
	x_new[329]=x[378]^x[374]^x[373]^x[372]^x[368]^x[367]^x[366]^x[363]^x[361]^x[357]^x[355]^x[351]^x[329]^x[276]^x[265]^x[255]^x[254]^x[249]^x[248]^x[245]^x[244]^x[243]^x[242]^x[239]^x[238]^x[237]^x[236]^x[234]^x[233]^x[231]^x[228]^x[227]^x[225]^x[214]^x[213]^x[212]^x[203]^x[201]^x[149]^x[148]^x[147]^x[139]^x[137]^x[128]^x[95]^x[94]^x[85]^x[84]^x[83]^x[82]^x[74]^x[73]^x[71]^x[41]^x[35];
	x_new[328]=x[373]^x[372]^x[371]^x[367]^x[366]^x[365]^x[362]^x[360]^x[356]^x[354]^x[350]^x[328]^x[275]^x[264]^x[254]^x[253]^x[248]^x[247]^x[244]^x[243]^x[242]^x[241]^x[238]^x[237]^x[236]^x[235]^x[233]^x[232]^x[230]^x[227]^x[226]^x[224]^x[213]^x[212]^x[211]^x[202]^x[200]^x[159]^x[148]^x[146]^x[136]^x[94]^x[93]^x[84]^x[83]^x[82]^x[81]^x[73]^x[72]^x[70]^x[40]^x[34];
	x_new[327]=x[372]^x[371]^x[370]^x[366]^x[365]^x[364]^x[361]^x[359]^x[355]^x[353]^x[349]^x[327]^x[274]^x[263]^x[253]^x[252]^x[247]^x[246]^x[243]^x[242]^x[241]^x[240]^x[237]^x[236]^x[235]^x[232]^x[231]^x[229]^x[226]^x[225]^x[212]^x[211]^x[210]^x[201]^x[199]^x[158]^x[147]^x[145]^x[135]^x[93]^x[92]^x[83]^x[82]^x[81]^x[80]^x[72]^x[71]^x[69]^x[39]^x[33];
	x_new[326]=x[371]^x[370]^x[369]^x[365]^x[364]^x[363]^x[360]^x[358]^x[354]^x[352]^x[348]^x[326]^x[273]^x[262]^x[252]^x[251]^x[246]^x[245]^x[242]^x[241]^x[240]^x[239]^x[236]^x[235]^x[234]^x[231]^x[230]^x[228]^x[225]^x[224]^x[211]^x[210]^x[209]^x[200]^x[198]^x[157]^x[146]^x[144]^x[134]^x[92]^x[91]^x[82]^x[81]^x[80]^x[79]^x[71]^x[70]^x[68]^x[38]^x[32];
	x_new[325]=x[374]^x[370]^x[369]^x[368]^x[359]^x[357]^x[352]^x[347]^x[325]^x[310]^x[288]^x[272]^x[261]^x[251]^x[250]^x[245]^x[244]^x[241]^x[240]^x[239]^x[238]^x[234]^x[233]^x[230]^x[229]^x[227]^x[210]^x[209]^x[208]^x[199]^x[197]^x[156]^x[145]^x[143]^x[106]^x[91]^x[90]^x[81]^x[80]^x[79]^x[78]^x[75]^x[70]^x[67]^x[64]^x[37];
	x_new[324]=x[369]^x[368]^x[367]^x[358]^x[356]^x[346]^x[324]^x[309]^x[298]^x[271]^x[260]^x[250]^x[249]^x[244]^x[243]^x[240]^x[239]^x[238]^x[237]^x[233]^x[232]^x[229]^x[228]^x[226]^x[209]^x[208]^x[207]^x[198]^x[196]^x[155]^x[144]^x[142]^x[132]^x[105]^x[90]^x[89]^x[80]^x[79]^x[78]^x[77]^x[74]^x[69]^x[66]^x[36];
	x_new[323]=x[368]^x[367]^x[366]^x[357]^x[355]^x[345]^x[323]^x[308]^x[297]^x[270]^x[259]^x[249]^x[248]^x[243]^x[242]^x[239]^x[238]^x[237]^x[236]^x[232]^x[231]^x[228]^x[227]^x[225]^x[208]^x[207]^x[206]^x[197]^x[195]^x[154]^x[143]^x[141]^x[131]^x[104]^x[89]^x[88]^x[79]^x[78]^x[77]^x[76]^x[73]^x[68]^x[65]^x[35];
	x_new[322]=x[367]^x[366]^x[365]^x[356]^x[354]^x[344]^x[322]^x[307]^x[296]^x[269]^x[258]^x[248]^x[247]^x[242]^x[241]^x[238]^x[237]^x[236]^x[235]^x[231]^x[230]^x[227]^x[226]^x[224]^x[207]^x[206]^x[205]^x[196]^x[194]^x[153]^x[142]^x[140]^x[130]^x[103]^x[88]^x[87]^x[78]^x[77]^x[76]^x[75]^x[72]^x[67]^x[64]^x[34];
	x_new[321]=x[366]^x[365]^x[364]^x[355]^x[353]^x[343]^x[321]^x[306]^x[295]^x[268]^x[257]^x[247]^x[246]^x[241]^x[240]^x[237]^x[236]^x[235]^x[230]^x[229]^x[226]^x[225]^x[206]^x[205]^x[204]^x[195]^x[193]^x[152]^x[141]^x[139]^x[129]^x[102]^x[87]^x[86]^x[77]^x[76]^x[75]^x[71]^x[66]^x[33];
	x_new[320]=x[365]^x[364]^x[363]^x[354]^x[352]^x[342]^x[320]^x[305]^x[294]^x[267]^x[256]^x[246]^x[240]^x[236]^x[235]^x[229]^x[225]^x[224]^x[205]^x[204]^x[203]^x[194]^x[192]^x[151]^x[140]^x[139]^x[101]^x[86]^x[76]^x[75]^x[70]^x[65]^x[32];
	x_new[319]=x[380]^x[369]^x[351]^x[347]^x[346]^x[345]^x[343]^x[342]^x[341]^x[337]^x[335]^x[331]^x[330]^x[326]^x[325]^x[324]^x[321]^x[319]^x[309]^x[299]^x[288]^x[282]^x[281]^x[272]^x[270]^x[261]^x[255]^x[254]^x[245]^x[243]^x[234]^x[221]^x[218]^x[215]^x[214]^x[212]^x[210]^x[208]^x[206]^x[204]^x[203]^x[202]^x[199]^x[197]^x[196]^x[193]^x[191]^x[183]^x[182]^x[181]^x[171]^x[170]^x[161]^x[145]^x[139]^x[117]^x[116]^x[115]^x[108]^x[107]^x[97]^x[96]^x[61]^x[58]^x[54]^x[50]^x[46]^x[43]^x[42]^x[40]^x[39]^x[31]^x[25]^x[19]^x[13];
	x_new[318]=x[379]^x[368]^x[350]^x[344]^x[342]^x[341]^x[340]^x[336]^x[335]^x[334]^x[330]^x[329]^x[325]^x[324]^x[323]^x[320]^x[319]^x[318]^x[308]^x[254]^x[253]^x[244]^x[242]^x[233]^x[222]^x[220]^x[216]^x[214]^x[213]^x[210]^x[209]^x[207]^x[204]^x[203]^x[202]^x[201]^x[199]^x[198]^x[196]^x[195]^x[193]^x[192]^x[190]^x[182]^x[181]^x[180]^x[170]^x[169]^x[160]^x[144]^x[138]^x[126]^x[114]^x[107]^x[106]^x[96]^x[62]^x[60]^x[53]^x[50]^x[49]^x[42]^x[41]^x[39]^x[38]^x[30]^x[24]^x[18]^x[12];
	x_new[317]=x[378]^x[367]^x[351]^x[349]^x[345]^x[343]^x[341]^x[340]^x[339]^x[335]^x[334]^x[333]^x[330]^x[329]^x[328]^x[324]^x[323]^x[322]^x[318]^x[317]^x[307]^x[253]^x[252]^x[243]^x[241]^x[232]^x[221]^x[219]^x[215]^x[213]^x[212]^x[209]^x[208]^x[206]^x[202]^x[201]^x[200]^x[198]^x[197]^x[195]^x[194]^x[191]^x[189]^x[181]^x[180]^x[179]^x[170]^x[169]^x[168]^x[143]^x[137]^x[127]^x[125]^x[115]^x[113]^x[105]^x[61]^x[59]^x[52]^x[49]^x[48]^x[41]^x[40]^x[38]^x[37]^x[29]^x[23]^x[17]^x[11];
	x_new[316]=x[377]^x[366]^x[350]^x[348]^x[344]^x[342]^x[340]^x[339]^x[338]^x[334]^x[333]^x[332]^x[329]^x[328]^x[327]^x[323]^x[322]^x[321]^x[317]^x[316]^x[306]^x[252]^x[251]^x[242]^x[240]^x[231]^x[220]^x[218]^x[214]^x[212]^x[211]^x[208]^x[207]^x[205]^x[201]^x[200]^x[199]^x[197]^x[196]^x[194]^x[193]^x[190]^x[188]^x[180]^x[179]^x[178]^x[169]^x[168]^x[167]^x[142]^x[136]^x[126]^x[124]^x[114]^x[112]^x[104]^x[60]^x[58]^x[51]^x[48]^x[47]^x[40]^x[39]^x[37]^x[36]^x[28]^x[22]^x[16]^x[10];
	x_new[315]=x[376]^x[365]^x[349]^x[347]^x[343]^x[341]^x[339]^x[338]^x[337]^x[333]^x[332]^x[331]^x[328]^x[327]^x[326]^x[322]^x[321]^x[320]^x[316]^x[315]^x[305]^x[251]^x[250]^x[241]^x[239]^x[230]^x[219]^x[217]^x[213]^x[211]^x[210]^x[207]^x[206]^x[204]^x[200]^x[199]^x[198]^x[196]^x[195]^x[193]^x[192]^x[189]^x[187]^x[179]^x[178]^x[177]^x[168]^x[167]^x[166]^x[141]^x[135]^x[125]^x[123]^x[113]^x[111]^x[103]^x[59]^x[57]^x[50]^x[47]^x[46]^x[39]^x[38]^x[36]^x[35]^x[27]^x[21]^x[15]^x[9];
	x_new[314]=x[375]^x[364]^x[351]^x[348]^x[346]^x[341]^x[340]^x[338]^x[337]^x[336]^x[332]^x[327]^x[326]^x[325]^x[321]^x[320]^x[315]^x[314]^x[304]^x[287]^x[286]^x[277]^x[276]^x[275]^x[267]^x[256]^x[250]^x[249]^x[240]^x[238]^x[229]^x[221]^x[218]^x[216]^x[213]^x[211]^x[210]^x[209]^x[206]^x[205]^x[203]^x[201]^x[198]^x[197]^x[195]^x[194]^x[192]^x[188]^x[186]^x[178]^x[177]^x[176]^x[167]^x[166]^x[165]^x[140]^x[134]^x[124]^x[112]^x[110]^x[102]^x[101]^x[95]^x[74]^x[58]^x[56]^x[53]^x[52]^x[51]^x[49]^x[47]^x[38]^x[37]^x[35]^x[34]^x[26]^x[20]^x[14]^x[8];
	x_new[313]=x[374]^x[363]^x[351]^x[350]^x[347]^x[345]^x[341]^x[340]^x[339]^x[337]^x[336]^x[335]^x[331]^x[326]^x[325]^x[324]^x[320]^x[314]^x[313]^x[303]^x[285]^x[276]^x[274]^x[249]^x[248]^x[239]^x[237]^x[228]^x[223]^x[220]^x[217]^x[215]^x[212]^x[210]^x[209]^x[208]^x[205]^x[204]^x[200]^x[197]^x[196]^x[194]^x[193]^x[187]^x[185]^x[177]^x[176]^x[175]^x[166]^x[165]^x[164]^x[139]^x[133]^x[123]^x[121]^x[111]^x[109]^x[101]^x[94]^x[73]^x[63]^x[55]^x[52]^x[50]^x[48]^x[46]^x[45]^x[42]^x[37]^x[34]^x[33]^x[25]^x[19]^x[13]^x[7];
	x_new[312]=x[373]^x[362]^x[351]^x[350]^x[349]^x[346]^x[344]^x[340]^x[339]^x[338]^x[336]^x[335]^x[334]^x[325]^x[324]^x[323]^x[313]^x[312]^x[302]^x[284]^x[275]^x[273]^x[248]^x[247]^x[238]^x[236]^x[227]^x[222]^x[219]^x[216]^x[214]^x[211]^x[209]^x[208]^x[207]^x[204]^x[203]^x[199]^x[196]^x[195]^x[193]^x[192]^x[186]^x[184]^x[176]^x[175]^x[174]^x[165]^x[164]^x[163]^x[138]^x[132]^x[122]^x[120]^x[110]^x[108]^x[100]^x[93]^x[72]^x[62]^x[54]^x[51]^x[49]^x[47]^x[45]^x[44]^x[41]^x[36]^x[33]^x[32]^x[24]^x[18]^x[12]^x[6];
	x_new[311]=x[372]^x[361]^x[350]^x[349]^x[348]^x[345]^x[343]^x[339]^x[338]^x[337]^x[335]^x[334]^x[333]^x[324]^x[323]^x[322]^x[312]^x[311]^x[301]^x[283]^x[274]^x[272]^x[247]^x[246]^x[237]^x[235]^x[226]^x[221]^x[218]^x[215]^x[210]^x[208]^x[206]^x[198]^x[196]^x[195]^x[194]^x[185]^x[183]^x[175]^x[174]^x[173]^x[164]^x[163]^x[162]^x[137]^x[131]^x[121]^x[119]^x[109]^x[107]^x[99]^x[92]^x[71]^x[61]^x[50]^x[48]^x[46]^x[44]^x[42]^x[40]^x[35]^x[23]^x[17]^x[11]^x[5];
	x_new[310]=x[371]^x[360]^x[349]^x[348]^x[347]^x[344]^x[342]^x[338]^x[337]^x[336]^x[334]^x[333]^x[332]^x[323]^x[322]^x[321]^x[311]^x[310]^x[300]^x[282]^x[273]^x[271]^x[246]^x[245]^x[236]^x[234]^x[225]^x[220]^x[217]^x[214]^x[209]^x[207]^x[205]^x[197]^x[195]^x[194]^x[193]^x[184]^x[182]^x[174]^x[173]^x[172]^x[163]^x[162]^x[161]^x[136]^x[130]^x[120]^x[118]^x[108]^x[106]^x[98]^x[91]^x[70]^x[60]^x[49]^x[47]^x[45]^x[43]^x[41]^x[39]^x[34]^x[22]^x[16]^x[10]^x[4];
	x_new[309]=x[370]^x[359]^x[348]^x[347]^x[346]^x[343]^x[341]^x[337]^x[336]^x[335]^x[333]^x[332]^x[331]^x[322]^x[321]^x[320]^x[310]^x[309]^x[299]^x[281]^x[272]^x[270]^x[245]^x[244]^x[235]^x[233]^x[224]^x[219]^x[216]^x[208]^x[207]^x[206]^x[204]^x[202]^x[194]^x[193]^x[192]^x[183]^x[181]^x[173]^x[172]^x[171]^x[162]^x[161]^x[160]^x[135]^x[129]^x[119]^x[117]^x[106]^x[105]^x[97]^x[96]^x[90]^x[69]^x[59]^x[53]^x[48]^x[46]^x[44]^x[40]^x[38]^x[33]^x[21]^x[15]^x[9]^x[3];
	x_new[308]=x[369]^x[358]^x[351]^x[347]^x[346]^x[345]^x[342]^x[340]^x[334]^x[332]^x[331]^x[325]^x[321]^x[320]^x[309]^x[308]^x[298]^x[282]^x[281]^x[270]^x[255]^x[244]^x[243]^x[232]^x[223]^x[222]^x[221]^x[218]^x[217]^x[216]^x[215]^x[212]^x[210]^x[206]^x[204]^x[203]^x[202]^x[196]^x[192]^x[191]^x[182]^x[180]^x[172]^x[171]^x[161]^x[160]^x[134]^x[128]^x[127]^x[126]^x[118]^x[106]^x[105]^x[104]^x[96]^x[63]^x[62]^x[61]^x[58]^x[50]^x[46]^x[43]^x[42]^x[40]^x[37]^x[32]^x[20]^x[14]^x[8]^x[2];
	x_new[307]=x[368]^x[357]^x[351]^x[350]^x[346]^x[345]^x[344]^x[341]^x[339]^x[335]^x[333]^x[331]^x[320]^x[308]^x[307]^x[297]^x[254]^x[243]^x[242]^x[231]^x[223]^x[222]^x[221]^x[220]^x[217]^x[216]^x[215]^x[214]^x[211]^x[209]^x[205]^x[203]^x[201]^x[195]^x[191]^x[190]^x[181]^x[179]^x[171]^x[160]^x[133]^x[127]^x[125]^x[117]^x[115]^x[106]^x[105]^x[104]^x[103]^x[63]^x[62]^x[61]^x[60]^x[51]^x[49]^x[41]^x[19]^x[13]^x[7]^x[1];
	x_new[306]=x[367]^x[356]^x[351]^x[350]^x[349]^x[345]^x[344]^x[343]^x[340]^x[338]^x[334]^x[332]^x[307]^x[306]^x[296]^x[253]^x[242]^x[241]^x[230]^x[222]^x[221]^x[220]^x[219]^x[216]^x[215]^x[214]^x[213]^x[210]^x[208]^x[204]^x[202]^x[200]^x[194]^x[191]^x[190]^x[189]^x[180]^x[178]^x[132]^x[126]^x[124]^x[116]^x[114]^x[105]^x[104]^x[103]^x[102]^x[62]^x[61]^x[60]^x[59]^x[50]^x[48]^x[40]^x[18]^x[12]^x[6]^x[0];
	x_new[305]=x[366]^x[355]^x[350]^x[349]^x[348]^x[344]^x[343]^x[342]^x[339]^x[337]^x[333]^x[331]^x[306]^x[305]^x[295]^x[278]^x[277]^x[266]^x[256]^x[252]^x[241]^x[240]^x[229]^x[221]^x[220]^x[219]^x[218]^x[215]^x[214]^x[213]^x[212]^x[209]^x[207]^x[202]^x[201]^x[199]^x[193]^x[192]^x[190]^x[189]^x[188]^x[179]^x[177]^x[131]^x[125]^x[123]^x[115]^x[113]^x[104]^x[103]^x[102]^x[101]^x[61]^x[60]^x[59]^x[58]^x[49]^x[47]^x[43]^x[42]^x[39]^x[37]^x[36]^x[32]^x[17]^x[11]^x[5];
	x_new[304]=x[365]^x[354]^x[349]^x[348]^x[347]^x[343]^x[342]^x[341]^x[338]^x[336]^x[332]^x[330]^x[305]^x[304]^x[294]^x[276]^x[265]^x[251]^x[240]^x[239]^x[228]^x[220]^x[219]^x[218]^x[217]^x[214]^x[213]^x[212]^x[211]^x[208]^x[206]^x[202]^x[201]^x[200]^x[198]^x[192]^x[189]^x[188]^x[187]^x[178]^x[176]^x[130]^x[124]^x[122]^x[114]^x[112]^x[103]^x[102]^x[101]^x[100]^x[60]^x[59]^x[58]^x[57]^x[48]^x[46]^x[41]^x[38]^x[35]^x[16]^x[10]^x[4];
	x_new[303]=x[364]^x[353]^x[348]^x[347]^x[346]^x[342]^x[341]^x[340]^x[337]^x[335]^x[330]^x[329]^x[320]^x[304]^x[303]^x[293]^x[277]^x[275]^x[266]^x[264]^x[250]^x[239]^x[238]^x[227]^x[219]^x[218]^x[217]^x[216]^x[213]^x[212]^x[211]^x[210]^x[207]^x[205]^x[202]^x[201]^x[200]^x[199]^x[197]^x[188]^x[187]^x[186]^x[177]^x[175]^x[129]^x[123]^x[121]^x[113]^x[111]^x[102]^x[101]^x[100]^x[99]^x[59]^x[58]^x[57]^x[56]^x[47]^x[45]^x[42]^x[40]^x[37]^x[36]^x[34]^x[15]^x[9]^x[3];
	x_new[302]=x[363]^x[352]^x[347]^x[346]^x[345]^x[341]^x[340]^x[339]^x[336]^x[334]^x[330]^x[329]^x[328]^x[303]^x[302]^x[292]^x[276]^x[274]^x[265]^x[263]^x[249]^x[238]^x[237]^x[226]^x[218]^x[217]^x[216]^x[215]^x[212]^x[211]^x[210]^x[209]^x[206]^x[204]^x[201]^x[200]^x[199]^x[198]^x[196]^x[187]^x[186]^x[185]^x[176]^x[174]^x[128]^x[122]^x[120]^x[112]^x[110]^x[101]^x[100]^x[99]^x[98]^x[58]^x[57]^x[56]^x[55]^x[46]^x[44]^x[41]^x[39]^x[36]^x[35]^x[33]^x[14]^x[8]^x[2];
	x_new[301]=x[346]^x[345]^x[344]^x[340]^x[339]^x[338]^x[335]^x[333]^x[329]^x[328]^x[327]^x[302]^x[301]^x[291]^x[275]^x[273]^x[264]^x[262]^x[248]^x[237]^x[236]^x[225]^x[217]^x[216]^x[215]^x[214]^x[211]^x[210]^x[209]^x[208]^x[205]^x[203]^x[200]^x[199]^x[198]^x[197]^x[195]^x[186]^x[185]^x[184]^x[175]^x[173]^x[121]^x[119]^x[111]^x[109]^x[100]^x[99]^x[98]^x[97]^x[57]^x[56]^x[55]^x[54]^x[45]^x[43]^x[40]^x[38]^x[35]^x[34]^x[32]^x[13]^x[7]^x[1];
	x_new[300]=x[345]^x[344]^x[343]^x[339]^x[338]^x[337]^x[334]^x[332]^x[328]^x[327]^x[326]^x[301]^x[300]^x[290]^x[274]^x[272]^x[263]^x[261]^x[247]^x[236]^x[235]^x[224]^x[216]^x[215]^x[214]^x[210]^x[209]^x[208]^x[204]^x[199]^x[198]^x[197]^x[194]^x[185]^x[184]^x[183]^x[174]^x[172]^x[120]^x[118]^x[110]^x[108]^x[99]^x[98]^x[97]^x[96]^x[56]^x[55]^x[54]^x[44]^x[39]^x[37]^x[34]^x[33]^x[12]^x[6]^x[0];
	x_new[299]=x[344]^x[343]^x[342]^x[338]^x[337]^x[336]^x[333]^x[331]^x[327]^x[326]^x[325]^x[300]^x[299]^x[289]^x[273]^x[272]^x[262]^x[261]^x[246]^x[235]^x[215]^x[214]^x[209]^x[208]^x[198]^x[197]^x[193]^x[192]^x[184]^x[183]^x[182]^x[173]^x[171]^x[119]^x[118]^x[109]^x[98]^x[97]^x[96]^x[55]^x[54]^x[38]^x[37]^x[33]^x[11]^x[5];
	x_new[298]=x[343]^x[342]^x[341]^x[337]^x[336]^x[335]^x[332]^x[330]^x[326]^x[325]^x[324]^x[299]^x[298]^x[288]^x[272]^x[261]^x[245]^x[234]^x[214]^x[213]^x[208]^x[207]^x[202]^x[197]^x[196]^x[192]^x[183]^x[182]^x[181]^x[172]^x[170]^x[118]^x[108]^x[106]^x[97]^x[96]^x[54]^x[53]^x[42]^x[37]^x[32]^x[10]^x[4];
	x_new[297]=x[346]^x[342]^x[341]^x[340]^x[336]^x[335]^x[334]^x[331]^x[329]^x[325]^x[323]^x[319]^x[297]^x[244]^x[233]^x[223]^x[222]^x[217]^x[216]^x[213]^x[212]^x[211]^x[210]^x[207]^x[206]^x[205]^x[204]^x[202]^x[201]^x[199]^x[196]^x[195]^x[193]^x[182]^x[181]^x[180]^x[171]^x[169]^x[117]^x[116]^x[115]^x[107]^x[105]^x[96]^x[63]^x[62]^x[53]^x[52]^x[51]^x[50]^x[42]^x[41]^x[39]^x[9]^x[3];
	x_new[296]=x[341]^x[340]^x[339]^x[335]^x[334]^x[333]^x[330]^x[328]^x[324]^x[322]^x[318]^x[296]^x[243]^x[232]^x[222]^x[221]^x[216]^x[215]^x[212]^x[211]^x[210]^x[209]^x[206]^x[205]^x[204]^x[203]^x[201]^x[200]^x[198]^x[195]^x[194]^x[192]^x[181]^x[180]^x[179]^x[170]^x[168]^x[127]^x[116]^x[114]^x[104]^x[62]^x[61]^x[52]^x[51]^x[50]^x[49]^x[41]^x[40]^x[38]^x[8]^x[2];
	x_new[295]=x[340]^x[339]^x[338]^x[334]^x[333]^x[332]^x[329]^x[327]^x[323]^x[321]^x[317]^x[295]^x[242]^x[231]^x[221]^x[220]^x[215]^x[214]^x[211]^x[210]^x[209]^x[208]^x[205]^x[204]^x[203]^x[200]^x[199]^x[197]^x[194]^x[193]^x[180]^x[179]^x[178]^x[169]^x[167]^x[126]^x[115]^x[113]^x[103]^x[61]^x[60]^x[51]^x[50]^x[49]^x[48]^x[40]^x[39]^x[37]^x[7]^x[1];
	x_new[294]=x[339]^x[338]^x[337]^x[333]^x[332]^x[331]^x[328]^x[326]^x[322]^x[320]^x[316]^x[294]^x[241]^x[230]^x[220]^x[219]^x[214]^x[213]^x[210]^x[209]^x[208]^x[207]^x[204]^x[203]^x[202]^x[199]^x[198]^x[196]^x[193]^x[192]^x[179]^x[178]^x[177]^x[168]^x[166]^x[125]^x[114]^x[112]^x[102]^x[60]^x[59]^x[50]^x[49]^x[48]^x[47]^x[39]^x[38]^x[36]^x[6]^x[0];
	x_new[293]=x[342]^x[338]^x[337]^x[336]^x[327]^x[325]^x[320]^x[315]^x[293]^x[278]^x[256]^x[240]^x[229]^x[219]^x[218]^x[213]^x[212]^x[209]^x[208]^x[207]^x[206]^x[202]^x[201]^x[198]^x[197]^x[195]^x[178]^x[177]^x[176]^x[167]^x[165]^x[124]^x[113]^x[111]^x[74]^x[59]^x[58]^x[49]^x[48]^x[47]^x[46]^x[43]^x[38]^x[35]^x[32]^x[5];
	x_new[292]=x[337]^x[336]^x[335]^x[326]^x[324]^x[314]^x[292]^x[277]^x[266]^x[239]^x[228]^x[218]^x[217]^x[212]^x[211]^x[208]^x[207]^x[206]^x[205]^x[201]^x[200]^x[197]^x[196]^x[194]^x[177]^x[176]^x[175]^x[166]^x[164]^x[123]^x[112]^x[110]^x[100]^x[73]^x[58]^x[57]^x[48]^x[47]^x[46]^x[45]^x[42]^x[37]^x[34]^x[4];
	x_new[291]=x[336]^x[335]^x[334]^x[325]^x[323]^x[313]^x[291]^x[276]^x[265]^x[238]^x[227]^x[217]^x[216]^x[211]^x[210]^x[207]^x[206]^x[205]^x[204]^x[200]^x[199]^x[196]^x[195]^x[193]^x[176]^x[175]^x[174]^x[165]^x[163]^x[122]^x[111]^x[109]^x[99]^x[72]^x[57]^x[56]^x[47]^x[46]^x[45]^x[44]^x[41]^x[36]^x[33]^x[3];
	x_new[290]=x[335]^x[334]^x[333]^x[324]^x[322]^x[312]^x[290]^x[275]^x[264]^x[237]^x[226]^x[216]^x[215]^x[210]^x[209]^x[206]^x[205]^x[204]^x[203]^x[199]^x[198]^x[195]^x[194]^x[192]^x[175]^x[174]^x[173]^x[164]^x[162]^x[121]^x[110]^x[108]^x[98]^x[71]^x[56]^x[55]^x[46]^x[45]^x[44]^x[43]^x[40]^x[35]^x[32]^x[2];
	x_new[289]=x[334]^x[333]^x[332]^x[323]^x[321]^x[311]^x[289]^x[274]^x[263]^x[236]^x[225]^x[215]^x[214]^x[209]^x[208]^x[205]^x[204]^x[203]^x[198]^x[197]^x[194]^x[193]^x[174]^x[173]^x[172]^x[163]^x[161]^x[120]^x[109]^x[107]^x[97]^x[70]^x[55]^x[54]^x[45]^x[44]^x[43]^x[39]^x[34]^x[1];
	x_new[288]=x[333]^x[332]^x[331]^x[322]^x[320]^x[310]^x[288]^x[273]^x[262]^x[235]^x[224]^x[214]^x[208]^x[204]^x[203]^x[197]^x[193]^x[192]^x[173]^x[172]^x[171]^x[162]^x[160]^x[119]^x[108]^x[107]^x[69]^x[54]^x[44]^x[43]^x[38]^x[33]^x[0];
	x_new[287]=x[383]^x[382]^x[377]^x[376]^x[373]^x[371]^x[367]^x[365]^x[362]^x[356]^x[348]^x[337]^x[319]^x[315]^x[314]^x[313]^x[311]^x[310]^x[309]^x[305]^x[303]^x[299]^x[298]^x[294]^x[293]^x[292]^x[289]^x[287]^x[277]^x[267]^x[256]^x[250]^x[249]^x[240]^x[238]^x[229]^x[223]^x[222]^x[213]^x[211]^x[202]^x[189]^x[186]^x[183]^x[182]^x[180]^x[178]^x[176]^x[174]^x[172]^x[171]^x[170]^x[167]^x[165]^x[164]^x[161]^x[151]^x[150]^x[149]^x[139]^x[138]^x[135]^x[129]^x[113]^x[107]^x[85]^x[84]^x[83]^x[76]^x[75]^x[65]^x[64]^x[29]^x[26]^x[22]^x[18]^x[14]^x[11]^x[10]^x[8]^x[7];
	x_new[286]=x[382]^x[381]^x[376]^x[375]^x[372]^x[370]^x[366]^x[364]^x[361]^x[355]^x[347]^x[336]^x[318]^x[312]^x[310]^x[309]^x[308]^x[304]^x[303]^x[302]^x[298]^x[297]^x[293]^x[292]^x[291]^x[288]^x[287]^x[286]^x[276]^x[222]^x[221]^x[212]^x[210]^x[201]^x[190]^x[188]^x[184]^x[182]^x[181]^x[178]^x[177]^x[175]^x[172]^x[171]^x[170]^x[169]^x[167]^x[166]^x[164]^x[163]^x[161]^x[160]^x[150]^x[149]^x[148]^x[138]^x[137]^x[134]^x[128]^x[112]^x[106]^x[94]^x[82]^x[75]^x[74]^x[64]^x[30]^x[28]^x[21]^x[18]^x[17]^x[10]^x[9]^x[7]^x[6];
	x_new[285]=x[381]^x[380]^x[375]^x[374]^x[371]^x[369]^x[365]^x[363]^x[360]^x[354]^x[346]^x[335]^x[319]^x[317]^x[313]^x[311]^x[309]^x[308]^x[307]^x[303]^x[302]^x[301]^x[298]^x[297]^x[296]^x[292]^x[291]^x[290]^x[286]^x[285]^x[275]^x[221]^x[220]^x[211]^x[209]^x[200]^x[189]^x[187]^x[183]^x[181]^x[180]^x[177]^x[176]^x[174]^x[170]^x[169]^x[168]^x[166]^x[165]^x[163]^x[162]^x[159]^x[149]^x[148]^x[147]^x[138]^x[137]^x[136]^x[133]^x[111]^x[105]^x[95]^x[93]^x[83]^x[81]^x[73]^x[29]^x[27]^x[20]^x[17]^x[16]^x[9]^x[8]^x[6]^x[5];
	x_new[284]=x[380]^x[379]^x[374]^x[373]^x[370]^x[368]^x[364]^x[362]^x[359]^x[353]^x[345]^x[334]^x[318]^x[316]^x[312]^x[310]^x[308]^x[307]^x[306]^x[302]^x[301]^x[300]^x[297]^x[296]^x[295]^x[291]^x[290]^x[289]^x[285]^x[284]^x[274]^x[220]^x[219]^x[210]^x[208]^x[199]^x[188]^x[186]^x[182]^x[180]^x[179]^x[176]^x[175]^x[173]^x[169]^x[168]^x[167]^x[165]^x[164]^x[162]^x[161]^x[158]^x[148]^x[147]^x[146]^x[137]^x[136]^x[135]^x[132]^x[110]^x[104]^x[94]^x[92]^x[82]^x[80]^x[72]^x[28]^x[26]^x[19]^x[16]^x[15]^x[8]^x[7]^x[5]^x[4];
	x_new[283]=x[379]^x[378]^x[373]^x[372]^x[369]^x[367]^x[363]^x[361]^x[358]^x[352]^x[344]^x[333]^x[317]^x[315]^x[311]^x[309]^x[307]^x[306]^x[305]^x[301]^x[300]^x[299]^x[296]^x[295]^x[294]^x[290]^x[289]^x[288]^x[284]^x[283]^x[273]^x[219]^x[218]^x[209]^x[207]^x[198]^x[187]^x[185]^x[181]^x[179]^x[178]^x[175]^x[174]^x[172]^x[168]^x[167]^x[166]^x[164]^x[163]^x[161]^x[160]^x[157]^x[147]^x[146]^x[145]^x[136]^x[135]^x[134]^x[131]^x[109]^x[103]^x[93]^x[91]^x[81]^x[79]^x[71]^x[27]^x[25]^x[18]^x[15]^x[14]^x[7]^x[6]^x[4]^x[3];
	x_new[282]=x[383]^x[378]^x[377]^x[372]^x[371]^x[368]^x[366]^x[360]^x[357]^x[343]^x[332]^x[319]^x[316]^x[314]^x[309]^x[308]^x[306]^x[305]^x[304]^x[300]^x[295]^x[294]^x[293]^x[289]^x[288]^x[283]^x[282]^x[272]^x[255]^x[254]^x[245]^x[244]^x[243]^x[235]^x[224]^x[218]^x[217]^x[208]^x[206]^x[197]^x[189]^x[186]^x[184]^x[181]^x[179]^x[178]^x[177]^x[174]^x[173]^x[171]^x[169]^x[166]^x[165]^x[163]^x[162]^x[160]^x[156]^x[146]^x[145]^x[144]^x[135]^x[134]^x[133]^x[130]^x[108]^x[102]^x[92]^x[80]^x[78]^x[70]^x[69]^x[63]^x[42]^x[26]^x[24]^x[21]^x[20]^x[19]^x[17]^x[15]^x[6]^x[5]^x[3]^x[2];
	x_new[281]=x[382]^x[377]^x[376]^x[371]^x[370]^x[367]^x[365]^x[359]^x[356]^x[342]^x[331]^x[319]^x[318]^x[315]^x[313]^x[309]^x[308]^x[307]^x[305]^x[304]^x[303]^x[299]^x[294]^x[293]^x[292]^x[288]^x[282]^x[281]^x[271]^x[253]^x[244]^x[242]^x[217]^x[216]^x[207]^x[205]^x[196]^x[191]^x[188]^x[185]^x[183]^x[180]^x[178]^x[177]^x[176]^x[173]^x[172]^x[168]^x[165]^x[164]^x[162]^x[161]^x[155]^x[145]^x[144]^x[143]^x[134]^x[133]^x[132]^x[129]^x[107]^x[101]^x[91]^x[89]^x[79]^x[77]^x[69]^x[62]^x[41]^x[31]^x[23]^x[20]^x[18]^x[16]^x[14]^x[13]^x[10]^x[5]^x[2]^x[1];
	x_new[280]=x[381]^x[376]^x[375]^x[370]^x[369]^x[366]^x[364]^x[358]^x[355]^x[341]^x[330]^x[319]^x[318]^x[317]^x[314]^x[312]^x[308]^x[307]^x[306]^x[304]^x[303]^x[302]^x[293]^x[292]^x[291]^x[281]^x[280]^x[270]^x[252]^x[243]^x[241]^x[216]^x[215]^x[206]^x[204]^x[195]^x[190]^x[187]^x[184]^x[182]^x[179]^x[177]^x[176]^x[175]^x[172]^x[171]^x[167]^x[164]^x[163]^x[161]^x[160]^x[154]^x[144]^x[143]^x[142]^x[133]^x[132]^x[131]^x[128]^x[106]^x[100]^x[90]^x[88]^x[78]^x[76]^x[68]^x[61]^x[40]^x[30]^x[22]^x[19]^x[17]^x[15]^x[13]^x[12]^x[9]^x[4]^x[1]^x[0];
	x_new[279]=x[380]^x[375]^x[374]^x[369]^x[368]^x[365]^x[363]^x[357]^x[354]^x[340]^x[329]^x[318]^x[317]^x[316]^x[313]^x[311]^x[307]^x[306]^x[305]^x[303]^x[302]^x[301]^x[292]^x[291]^x[290]^x[280]^x[279]^x[269]^x[251]^x[242]^x[240]^x[215]^x[214]^x[205]^x[203]^x[194]^x[189]^x[186]^x[183]^x[178]^x[176]^x[174]^x[166]^x[164]^x[163]^x[162]^x[153]^x[143]^x[142]^x[141]^x[132]^x[131]^x[130]^x[105]^x[99]^x[89]^x[87]^x[77]^x[75]^x[67]^x[60]^x[39]^x[29]^x[18]^x[16]^x[14]^x[12]^x[10]^x[8]^x[3];
	x_new[278]=x[379]^x[374]^x[373]^x[368]^x[367]^x[364]^x[362]^x[356]^x[353]^x[339]^x[328]^x[317]^x[316]^x[315]^x[312]^x[310]^x[306]^x[305]^x[304]^x[302]^x[301]^x[300]^x[291]^x[290]^x[289]^x[279]^x[278]^x[268]^x[250]^x[241]^x[239]^x[214]^x[213]^x[204]^x[202]^x[193]^x[188]^x[185]^x[182]^x[177]^x[175]^x[173]^x[165]^x[163]^x[162]^x[161]^x[152]^x[142]^x[141]^x[140]^x[131]^x[130]^x[129]^x[104]^x[98]^x[88]^x[86]^x[76]^x[74]^x[66]^x[59]^x[38]^x[28]^x[17]^x[15]^x[13]^x[11]^x[9]^x[7]^x[2];
	x_new[277]=x[378]^x[373]^x[372]^x[367]^x[366]^x[363]^x[361]^x[355]^x[352]^x[338]^x[327]^x[316]^x[315]^x[314]^x[311]^x[309]^x[305]^x[304]^x[303]^x[301]^x[300]^x[299]^x[290]^x[289]^x[288]^x[278]^x[277]^x[267]^x[249]^x[240]^x[238]^x[213]^x[212]^x[203]^x[201]^x[192]^x[187]^x[184]^x[176]^x[175]^x[174]^x[172]^x[170]^x[162]^x[161]^x[160]^x[151]^x[141]^x[140]^x[139]^x[130]^x[129]^x[128]^x[103]^x[97]^x[87]^x[85]^x[74]^x[73]^x[65]^x[64]^x[58]^x[37]^x[27]^x[21]^x[16]^x[14]^x[12]^x[8]^x[6]^x[1];
	x_new[276]=x[383]^x[377]^x[372]^x[371]^x[366]^x[365]^x[360]^x[354]^x[337]^x[326]^x[319]^x[315]^x[314]^x[313]^x[310]^x[308]^x[302]^x[300]^x[299]^x[293]^x[289]^x[288]^x[277]^x[276]^x[266]^x[250]^x[249]^x[238]^x[223]^x[212]^x[211]^x[200]^x[191]^x[190]^x[189]^x[186]^x[185]^x[184]^x[183]^x[180]^x[178]^x[174]^x[172]^x[171]^x[170]^x[164]^x[160]^x[159]^x[150]^x[140]^x[139]^x[129]^x[128]^x[102]^x[96]^x[95]^x[94]^x[86]^x[74]^x[73]^x[72]^x[64]^x[31]^x[30]^x[29]^x[26]^x[18]^x[14]^x[11]^x[10]^x[8]^x[5]^x[0];
	x_new[275]=x[382]^x[376]^x[371]^x[370]^x[365]^x[364]^x[359]^x[353]^x[336]^x[325]^x[319]^x[318]^x[314]^x[313]^x[312]^x[309]^x[307]^x[303]^x[301]^x[299]^x[288]^x[276]^x[275]^x[265]^x[222]^x[211]^x[210]^x[199]^x[191]^x[190]^x[189]^x[188]^x[185]^x[184]^x[183]^x[182]^x[179]^x[177]^x[173]^x[171]^x[169]^x[163]^x[159]^x[158]^x[149]^x[139]^x[128]^x[101]^x[95]^x[93]^x[85]^x[83]^x[74]^x[73]^x[72]^x[71]^x[31]^x[30]^x[29]^x[28]^x[19]^x[17]^x[9];
	x_new[274]=x[381]^x[375]^x[370]^x[369]^x[364]^x[363]^x[358]^x[352]^x[335]^x[324]^x[319]^x[318]^x[317]^x[313]^x[312]^x[311]^x[308]^x[306]^x[302]^x[300]^x[275]^x[274]^x[264]^x[221]^x[210]^x[209]^x[198]^x[190]^x[189]^x[188]^x[187]^x[184]^x[183]^x[182]^x[181]^x[178]^x[176]^x[172]^x[170]^x[168]^x[162]^x[159]^x[158]^x[157]^x[148]^x[100]^x[94]^x[92]^x[84]^x[82]^x[73]^x[72]^x[71]^x[70]^x[30]^x[29]^x[28]^x[27]^x[18]^x[16]^x[8];
	x_new[273]=x[380]^x[374]^x[369]^x[368]^x[363]^x[357]^x[334]^x[323]^x[318]^x[317]^x[316]^x[312]^x[311]^x[310]^x[307]^x[305]^x[301]^x[299]^x[274]^x[273]^x[263]^x[246]^x[245]^x[234]^x[224]^x[220]^x[209]^x[208]^x[197]^x[189]^x[188]^x[187]^x[186]^x[183]^x[182]^x[181]^x[180]^x[177]^x[175]^x[170]^x[169]^x[167]^x[161]^x[160]^x[158]^x[157]^x[156]^x[147]^x[99]^x[93]^x[91]^x[83]^x[81]^x[72]^x[71]^x[70]^x[69]^x[29]^x[28]^x[27]^x[26]^x[17]^x[15]^x[11]^x[10]^x[7]^x[5]^x[4]^x[0];
	x_new[272]=x[379]^x[373]^x[368]^x[367]^x[362]^x[356]^x[333]^x[322]^x[317]^x[316]^x[315]^x[311]^x[310]^x[309]^x[306]^x[304]^x[300]^x[298]^x[273]^x[272]^x[262]^x[244]^x[233]^x[219]^x[208]^x[207]^x[196]^x[188]^x[187]^x[186]^x[185]^x[182]^x[181]^x[180]^x[179]^x[176]^x[174]^x[170]^x[169]^x[168]^x[166]^x[160]^x[157]^x[156]^x[155]^x[146]^x[98]^x[92]^x[90]^x[82]^x[80]^x[71]^x[70]^x[69]^x[68]^x[28]^x[27]^x[26]^x[25]^x[16]^x[14]^x[9]^x[6]^x[3];
	x_new[271]=x[378]^x[372]^x[367]^x[366]^x[361]^x[355]^x[332]^x[321]^x[316]^x[315]^x[314]^x[310]^x[309]^x[308]^x[305]^x[303]^x[298]^x[297]^x[288]^x[272]^x[271]^x[261]^x[245]^x[243]^x[234]^x[232]^x[218]^x[207]^x[206]^x[195]^x[187]^x[186]^x[185]^x[184]^x[181]^x[180]^x[179]^x[178]^x[175]^x[173]^x[170]^x[169]^x[168]^x[167]^x[165]^x[156]^x[155]^x[154]^x[145]^x[97]^x[91]^x[89]^x[81]^x[79]^x[70]^x[69]^x[68]^x[67]^x[27]^x[26]^x[25]^x[24]^x[15]^x[13]^x[10]^x[8]^x[5]^x[4]^x[2];
	x_new[270]=x[377]^x[371]^x[366]^x[365]^x[360]^x[354]^x[331]^x[320]^x[315]^x[314]^x[313]^x[309]^x[308]^x[307]^x[304]^x[302]^x[298]^x[297]^x[296]^x[271]^x[270]^x[260]^x[244]^x[242]^x[233]^x[231]^x[217]^x[206]^x[205]^x[194]^x[186]^x[185]^x[184]^x[183]^x[180]^x[179]^x[178]^x[177]^x[174]^x[172]^x[169]^x[168]^x[167]^x[166]^x[164]^x[155]^x[154]^x[153]^x[144]^x[96]^x[90]^x[88]^x[80]^x[78]^x[69]^x[68]^x[67]^x[66]^x[26]^x[25]^x[24]^x[23]^x[14]^x[12]^x[9]^x[7]^x[4]^x[3]^x[1];
	x_new[269]=x[376]^x[370]^x[365]^x[364]^x[359]^x[353]^x[314]^x[313]^x[312]^x[308]^x[307]^x[306]^x[303]^x[301]^x[297]^x[296]^x[295]^x[270]^x[269]^x[259]^x[243]^x[241]^x[232]^x[230]^x[216]^x[205]^x[204]^x[193]^x[185]^x[184]^x[183]^x[182]^x[179]^x[178]^x[177]^x[176]^x[173]^x[171]^x[168]^x[167]^x[166]^x[165]^x[163]^x[154]^x[153]^x[152]^x[143]^x[89]^x[87]^x[79]^x[77]^x[68]^x[67]^x[66]^x[65]^x[25]^x[24]^x[23]^x[22]^x[13]^x[11]^x[8]^x[6]^x[3]^x[2]^x[0];
	x_new[268]=x[375]^x[369]^x[364]^x[363]^x[358]^x[352]^x[313]^x[312]^x[311]^x[307]^x[306]^x[305]^x[302]^x[300]^x[296]^x[295]^x[294]^x[269]^x[268]^x[258]^x[242]^x[240]^x[231]^x[229]^x[215]^x[204]^x[203]^x[192]^x[184]^x[183]^x[182]^x[178]^x[177]^x[176]^x[172]^x[167]^x[166]^x[165]^x[162]^x[153]^x[152]^x[151]^x[142]^x[88]^x[86]^x[78]^x[76]^x[67]^x[66]^x[65]^x[64]^x[24]^x[23]^x[22]^x[12]^x[7]^x[5]^x[2]^x[1];
	x_new[267]=x[374]^x[368]^x[363]^x[357]^x[312]^x[311]^x[310]^x[306]^x[305]^x[304]^x[301]^x[299]^x[295]^x[294]^x[293]^x[268]^x[267]^x[257]^x[241]^x[240]^x[230]^x[229]^x[214]^x[203]^x[183]^x[182]^x[177]^x[176]^x[166]^x[165]^x[161]^x[160]^x[152]^x[151]^x[150]^x[141]^x[87]^x[86]^x[77]^x[66]^x[65]^x[64]^x[23]^x[22]^x[6]^x[5]^x[1];
	x_new[266]=x[373]^x[367]^x[362]^x[356]^x[311]^x[310]^x[309]^x[305]^x[304]^x[303]^x[300]^x[298]^x[294]^x[293]^x[292]^x[267]^x[266]^x[256]^x[240]^x[229]^x[213]^x[202]^x[182]^x[181]^x[176]^x[175]^x[170]^x[165]^x[164]^x[160]^x[151]^x[150]^x[149]^x[140]^x[86]^x[76]^x[74]^x[65]^x[64]^x[22]^x[21]^x[10]^x[5]^x[0];
	x_new[265]=x[372]^x[366]^x[361]^x[355]^x[314]^x[310]^x[309]^x[308]^x[304]^x[303]^x[302]^x[299]^x[297]^x[293]^x[291]^x[287]^x[265]^x[212]^x[201]^x[191]^x[190]^x[185]^x[184]^x[181]^x[180]^x[179]^x[178]^x[175]^x[174]^x[173]^x[172]^x[170]^x[169]^x[167]^x[164]^x[163]^x[161]^x[150]^x[149]^x[148]^x[139]^x[85]^x[84]^x[83]^x[75]^x[73]^x[64]^x[31]^x[30]^x[21]^x[20]^x[19]^x[18]^x[10]^x[9]^x[7];
	x_new[264]=x[371]^x[365]^x[360]^x[354]^x[309]^x[308]^x[307]^x[303]^x[302]^x[301]^x[298]^x[296]^x[292]^x[290]^x[286]^x[264]^x[211]^x[200]^x[190]^x[189]^x[184]^x[183]^x[180]^x[179]^x[178]^x[177]^x[174]^x[173]^x[172]^x[171]^x[169]^x[168]^x[166]^x[163]^x[162]^x[160]^x[149]^x[148]^x[147]^x[138]^x[95]^x[84]^x[82]^x[72]^x[30]^x[29]^x[20]^x[19]^x[18]^x[17]^x[9]^x[8]^x[6];
	x_new[263]=x[370]^x[364]^x[359]^x[353]^x[308]^x[307]^x[306]^x[302]^x[301]^x[300]^x[297]^x[295]^x[291]^x[289]^x[285]^x[263]^x[210]^x[199]^x[189]^x[188]^x[183]^x[182]^x[179]^x[178]^x[177]^x[176]^x[173]^x[172]^x[171]^x[168]^x[167]^x[165]^x[162]^x[161]^x[148]^x[147]^x[146]^x[137]^x[94]^x[83]^x[81]^x[71]^x[29]^x[28]^x[19]^x[18]^x[17]^x[16]^x[8]^x[7]^x[5];
	x_new[262]=x[369]^x[363]^x[358]^x[352]^x[307]^x[306]^x[305]^x[301]^x[300]^x[299]^x[296]^x[294]^x[290]^x[288]^x[284]^x[262]^x[209]^x[198]^x[188]^x[187]^x[182]^x[181]^x[178]^x[177]^x[176]^x[175]^x[172]^x[171]^x[170]^x[167]^x[166]^x[164]^x[161]^x[160]^x[147]^x[146]^x[145]^x[136]^x[93]^x[82]^x[80]^x[70]^x[28]^x[27]^x[18]^x[17]^x[16]^x[15]^x[7]^x[6]^x[4];
	x_new[261]=x[368]^x[357]^x[310]^x[306]^x[305]^x[304]^x[295]^x[293]^x[288]^x[283]^x[261]^x[246]^x[224]^x[208]^x[197]^x[187]^x[186]^x[181]^x[180]^x[177]^x[176]^x[175]^x[174]^x[170]^x[169]^x[166]^x[165]^x[163]^x[146]^x[145]^x[144]^x[135]^x[92]^x[81]^x[79]^x[42]^x[27]^x[26]^x[17]^x[16]^x[15]^x[14]^x[11]^x[6]^x[3]^x[0];
	x_new[260]=x[367]^x[356]^x[305]^x[304]^x[303]^x[294]^x[292]^x[282]^x[260]^x[245]^x[234]^x[207]^x[196]^x[186]^x[185]^x[180]^x[179]^x[176]^x[175]^x[174]^x[173]^x[169]^x[168]^x[165]^x[164]^x[162]^x[145]^x[144]^x[143]^x[134]^x[91]^x[80]^x[78]^x[68]^x[41]^x[26]^x[25]^x[16]^x[15]^x[14]^x[13]^x[10]^x[5]^x[2];
	x_new[259]=x[366]^x[355]^x[304]^x[303]^x[302]^x[293]^x[291]^x[281]^x[259]^x[244]^x[233]^x[206]^x[195]^x[185]^x[184]^x[179]^x[178]^x[175]^x[174]^x[173]^x[172]^x[168]^x[167]^x[164]^x[163]^x[161]^x[144]^x[143]^x[142]^x[133]^x[90]^x[79]^x[77]^x[67]^x[40]^x[25]^x[24]^x[15]^x[14]^x[13]^x[12]^x[9]^x[4]^x[1];
	x_new[258]=x[365]^x[354]^x[303]^x[302]^x[301]^x[292]^x[290]^x[280]^x[258]^x[243]^x[232]^x[205]^x[194]^x[184]^x[183]^x[178]^x[177]^x[174]^x[173]^x[172]^x[171]^x[167]^x[166]^x[163]^x[162]^x[160]^x[143]^x[142]^x[141]^x[132]^x[89]^x[78]^x[76]^x[66]^x[39]^x[24]^x[23]^x[14]^x[13]^x[12]^x[11]^x[8]^x[3]^x[0];
	x_new[257]=x[364]^x[353]^x[302]^x[301]^x[300]^x[291]^x[289]^x[279]^x[257]^x[242]^x[231]^x[204]^x[193]^x[183]^x[182]^x[177]^x[176]^x[173]^x[172]^x[171]^x[166]^x[165]^x[162]^x[161]^x[142]^x[141]^x[140]^x[131]^x[88]^x[77]^x[75]^x[65]^x[38]^x[23]^x[22]^x[13]^x[12]^x[11]^x[7]^x[2];
	x_new[256]=x[363]^x[352]^x[301]^x[300]^x[299]^x[290]^x[288]^x[278]^x[256]^x[241]^x[230]^x[203]^x[192]^x[182]^x[176]^x[172]^x[171]^x[165]^x[161]^x[160]^x[141]^x[140]^x[139]^x[130]^x[87]^x[76]^x[75]^x[37]^x[22]^x[12]^x[11]^x[6]^x[1];
	x_new[255]=x[378]^x[377]^x[373]^x[368]^x[366]^x[364]^x[363]^x[362]^x[359]^x[357]^x[353]^x[351]^x[350]^x[345]^x[344]^x[341]^x[339]^x[335]^x[333]^x[330]^x[324]^x[316]^x[305]^x[287]^x[283]^x[282]^x[281]^x[279]^x[278]^x[277]^x[273]^x[271]^x[267]^x[266]^x[262]^x[261]^x[260]^x[257]^x[255]^x[245]^x[235]^x[224]^x[218]^x[217]^x[208]^x[206]^x[197]^x[191]^x[190]^x[181]^x[179]^x[170]^x[130]^x[119]^x[118]^x[117]^x[107]^x[106]^x[103]^x[97]^x[81]^x[75]^x[53]^x[52]^x[51]^x[44]^x[43]^x[33]^x[32];
	x_new[254]=x[382]^x[381]^x[370]^x[363]^x[362]^x[358]^x[352]^x[350]^x[349]^x[344]^x[343]^x[340]^x[338]^x[334]^x[332]^x[329]^x[323]^x[315]^x[304]^x[286]^x[280]^x[278]^x[277]^x[276]^x[272]^x[271]^x[270]^x[266]^x[265]^x[261]^x[260]^x[259]^x[256]^x[255]^x[254]^x[244]^x[190]^x[189]^x[180]^x[178]^x[169]^x[118]^x[117]^x[116]^x[106]^x[105]^x[102]^x[96]^x[80]^x[74]^x[62]^x[50]^x[43]^x[42]^x[32];
	x_new[253]=x[383]^x[381]^x[380]^x[369]^x[361]^x[357]^x[349]^x[348]^x[343]^x[342]^x[339]^x[337]^x[333]^x[331]^x[328]^x[322]^x[314]^x[303]^x[287]^x[285]^x[281]^x[279]^x[277]^x[276]^x[275]^x[271]^x[270]^x[269]^x[266]^x[265]^x[264]^x[260]^x[259]^x[258]^x[254]^x[253]^x[243]^x[189]^x[188]^x[179]^x[177]^x[168]^x[139]^x[128]^x[127]^x[117]^x[116]^x[115]^x[106]^x[105]^x[104]^x[101]^x[79]^x[73]^x[63]^x[61]^x[51]^x[49]^x[41];
	x_new[252]=x[382]^x[380]^x[379]^x[368]^x[360]^x[356]^x[348]^x[347]^x[342]^x[341]^x[338]^x[336]^x[332]^x[330]^x[327]^x[321]^x[313]^x[302]^x[286]^x[284]^x[280]^x[278]^x[276]^x[275]^x[274]^x[270]^x[269]^x[268]^x[265]^x[264]^x[263]^x[259]^x[258]^x[257]^x[253]^x[252]^x[242]^x[188]^x[187]^x[178]^x[176]^x[167]^x[138]^x[126]^x[116]^x[115]^x[114]^x[105]^x[104]^x[103]^x[100]^x[78]^x[72]^x[62]^x[60]^x[50]^x[48]^x[40];
	x_new[251]=x[381]^x[379]^x[378]^x[367]^x[359]^x[355]^x[347]^x[346]^x[341]^x[340]^x[337]^x[335]^x[331]^x[329]^x[326]^x[320]^x[312]^x[301]^x[285]^x[283]^x[279]^x[277]^x[275]^x[274]^x[273]^x[269]^x[268]^x[267]^x[264]^x[263]^x[262]^x[258]^x[257]^x[256]^x[252]^x[251]^x[241]^x[187]^x[186]^x[177]^x[175]^x[166]^x[137]^x[125]^x[115]^x[114]^x[113]^x[104]^x[103]^x[102]^x[99]^x[77]^x[71]^x[61]^x[59]^x[49]^x[47]^x[39];
	x_new[250]=x[383]^x[382]^x[380]^x[376]^x[373]^x[372]^x[371]^x[367]^x[365]^x[363]^x[358]^x[354]^x[352]^x[351]^x[346]^x[345]^x[340]^x[339]^x[336]^x[334]^x[328]^x[325]^x[311]^x[300]^x[287]^x[284]^x[282]^x[277]^x[276]^x[274]^x[273]^x[272]^x[268]^x[263]^x[262]^x[261]^x[257]^x[256]^x[251]^x[250]^x[240]^x[223]^x[222]^x[213]^x[212]^x[211]^x[203]^x[192]^x[186]^x[185]^x[176]^x[174]^x[165]^x[157]^x[124]^x[114]^x[113]^x[112]^x[103]^x[102]^x[101]^x[98]^x[76]^x[70]^x[60]^x[48]^x[46]^x[38]^x[37]^x[31]^x[10];
	x_new[249]=x[381]^x[379]^x[377]^x[376]^x[375]^x[372]^x[370]^x[366]^x[365]^x[364]^x[357]^x[353]^x[350]^x[345]^x[344]^x[339]^x[338]^x[335]^x[333]^x[327]^x[324]^x[310]^x[299]^x[287]^x[286]^x[283]^x[281]^x[277]^x[276]^x[275]^x[273]^x[272]^x[271]^x[267]^x[262]^x[261]^x[260]^x[256]^x[250]^x[249]^x[239]^x[221]^x[212]^x[210]^x[185]^x[184]^x[175]^x[173]^x[164]^x[156]^x[135]^x[123]^x[113]^x[112]^x[111]^x[102]^x[101]^x[100]^x[97]^x[75]^x[69]^x[59]^x[57]^x[47]^x[45]^x[37]^x[30]^x[9];
	x_new[248]=x[380]^x[378]^x[376]^x[375]^x[374]^x[371]^x[369]^x[365]^x[364]^x[363]^x[356]^x[352]^x[349]^x[344]^x[343]^x[338]^x[337]^x[334]^x[332]^x[326]^x[323]^x[309]^x[298]^x[287]^x[286]^x[285]^x[282]^x[280]^x[276]^x[275]^x[274]^x[272]^x[271]^x[270]^x[261]^x[260]^x[259]^x[249]^x[248]^x[238]^x[220]^x[211]^x[209]^x[184]^x[183]^x[174]^x[172]^x[163]^x[155]^x[134]^x[122]^x[112]^x[111]^x[110]^x[101]^x[100]^x[99]^x[96]^x[74]^x[68]^x[58]^x[56]^x[46]^x[44]^x[36]^x[29]^x[8];
	x_new[247]=x[379]^x[377]^x[375]^x[373]^x[370]^x[368]^x[364]^x[362]^x[355]^x[348]^x[343]^x[342]^x[337]^x[336]^x[333]^x[331]^x[325]^x[322]^x[308]^x[297]^x[286]^x[285]^x[284]^x[281]^x[279]^x[275]^x[274]^x[273]^x[271]^x[270]^x[269]^x[260]^x[259]^x[258]^x[248]^x[247]^x[237]^x[219]^x[210]^x[208]^x[183]^x[182]^x[173]^x[171]^x[162]^x[154]^x[121]^x[111]^x[110]^x[109]^x[100]^x[99]^x[98]^x[73]^x[67]^x[57]^x[55]^x[45]^x[43]^x[35]^x[28]^x[7];
	x_new[246]=x[378]^x[376]^x[374]^x[372]^x[369]^x[367]^x[363]^x[361]^x[354]^x[347]^x[342]^x[341]^x[336]^x[335]^x[332]^x[330]^x[324]^x[321]^x[307]^x[296]^x[285]^x[284]^x[283]^x[280]^x[278]^x[274]^x[273]^x[272]^x[270]^x[269]^x[268]^x[259]^x[258]^x[257]^x[247]^x[246]^x[236]^x[218]^x[209]^x[207]^x[182]^x[181]^x[172]^x[170]^x[161]^x[153]^x[120]^x[110]^x[109]^x[108]^x[99]^x[98]^x[97]^x[72]^x[66]^x[56]^x[54]^x[44]^x[42]^x[34]^x[27]^x[6];
	x_new[245]=x[377]^x[375]^x[373]^x[371]^x[368]^x[366]^x[363]^x[360]^x[353]^x[352]^x[346]^x[341]^x[340]^x[335]^x[334]^x[331]^x[329]^x[323]^x[320]^x[306]^x[295]^x[284]^x[283]^x[282]^x[279]^x[277]^x[273]^x[272]^x[271]^x[269]^x[268]^x[267]^x[258]^x[257]^x[256]^x[246]^x[245]^x[235]^x[217]^x[208]^x[206]^x[181]^x[180]^x[171]^x[169]^x[160]^x[152]^x[119]^x[109]^x[108]^x[107]^x[98]^x[97]^x[96]^x[71]^x[65]^x[55]^x[53]^x[42]^x[41]^x[33]^x[32]^x[26]^x[5];
	x_new[244]=x[383]^x[382]^x[378]^x[377]^x[374]^x[372]^x[370]^x[366]^x[361]^x[352]^x[351]^x[345]^x[340]^x[339]^x[334]^x[333]^x[328]^x[322]^x[305]^x[294]^x[287]^x[283]^x[282]^x[281]^x[278]^x[276]^x[270]^x[268]^x[267]^x[261]^x[257]^x[256]^x[245]^x[244]^x[234]^x[218]^x[217]^x[206]^x[191]^x[180]^x[179]^x[168]^x[130]^x[127]^x[118]^x[108]^x[107]^x[97]^x[96]^x[70]^x[64]^x[63]^x[62]^x[54]^x[42]^x[41]^x[40]^x[32];
	x_new[243]=x[383]^x[381]^x[373]^x[370]^x[369]^x[362]^x[360]^x[359]^x[350]^x[344]^x[339]^x[338]^x[333]^x[332]^x[327]^x[321]^x[304]^x[293]^x[287]^x[286]^x[282]^x[281]^x[280]^x[277]^x[275]^x[271]^x[269]^x[267]^x[256]^x[244]^x[243]^x[233]^x[190]^x[179]^x[178]^x[167]^x[127]^x[126]^x[117]^x[107]^x[96]^x[69]^x[63]^x[61]^x[53]^x[51]^x[42]^x[41]^x[40]^x[39];
	x_new[242]=x[382]^x[380]^x[372]^x[369]^x[368]^x[361]^x[359]^x[358]^x[349]^x[343]^x[338]^x[337]^x[332]^x[331]^x[326]^x[320]^x[303]^x[292]^x[287]^x[286]^x[285]^x[281]^x[280]^x[279]^x[276]^x[274]^x[270]^x[268]^x[243]^x[242]^x[232]^x[189]^x[178]^x[177]^x[166]^x[127]^x[126]^x[125]^x[116]^x[68]^x[62]^x[60]^x[52]^x[50]^x[41]^x[40]^x[39]^x[38];
	x_new[241]=x[381]^x[379]^x[374]^x[373]^x[371]^x[362]^x[360]^x[358]^x[356]^x[352]^x[348]^x[342]^x[337]^x[336]^x[331]^x[325]^x[302]^x[291]^x[286]^x[285]^x[284]^x[280]^x[279]^x[278]^x[275]^x[273]^x[269]^x[267]^x[242]^x[241]^x[231]^x[214]^x[213]^x[202]^x[192]^x[188]^x[177]^x[176]^x[165]^x[126]^x[125]^x[124]^x[115]^x[67]^x[61]^x[59]^x[51]^x[49]^x[40]^x[39]^x[38]^x[37];
	x_new[240]=x[380]^x[378]^x[372]^x[370]^x[367]^x[361]^x[359]^x[357]^x[356]^x[355]^x[347]^x[341]^x[336]^x[335]^x[330]^x[324]^x[301]^x[290]^x[285]^x[284]^x[283]^x[279]^x[278]^x[277]^x[274]^x[272]^x[268]^x[266]^x[241]^x[240]^x[230]^x[212]^x[201]^x[187]^x[176]^x[175]^x[164]^x[125]^x[124]^x[123]^x[114]^x[66]^x[60]^x[58]^x[50]^x[48]^x[39]^x[38]^x[37]^x[36];
	x_new[239]=x[379]^x[377]^x[373]^x[371]^x[369]^x[367]^x[366]^x[362]^x[360]^x[358]^x[355]^x[354]^x[346]^x[340]^x[335]^x[334]^x[329]^x[323]^x[300]^x[289]^x[284]^x[283]^x[282]^x[278]^x[277]^x[276]^x[273]^x[271]^x[266]^x[265]^x[256]^x[240]^x[239]^x[229]^x[213]^x[211]^x[202]^x[200]^x[186]^x[175]^x[174]^x[163]^x[124]^x[123]^x[122]^x[113]^x[65]^x[59]^x[57]^x[49]^x[47]^x[38]^x[37]^x[36]^x[35];
	x_new[238]=x[378]^x[376]^x[372]^x[370]^x[368]^x[366]^x[365]^x[361]^x[359]^x[357]^x[354]^x[353]^x[345]^x[339]^x[334]^x[333]^x[328]^x[322]^x[299]^x[288]^x[283]^x[282]^x[281]^x[277]^x[276]^x[275]^x[272]^x[270]^x[266]^x[265]^x[264]^x[239]^x[238]^x[228]^x[212]^x[210]^x[201]^x[199]^x[185]^x[174]^x[173]^x[162]^x[123]^x[122]^x[121]^x[112]^x[64]^x[58]^x[56]^x[48]^x[46]^x[37]^x[36]^x[35]^x[34];
	x_new[237]=x[377]^x[375]^x[371]^x[369]^x[367]^x[365]^x[364]^x[360]^x[358]^x[356]^x[353]^x[352]^x[344]^x[338]^x[333]^x[332]^x[327]^x[321]^x[282]^x[281]^x[280]^x[276]^x[275]^x[274]^x[271]^x[269]^x[265]^x[264]^x[263]^x[238]^x[237]^x[227]^x[211]^x[209]^x[200]^x[198]^x[184]^x[173]^x[172]^x[161]^x[122]^x[121]^x[120]^x[111]^x[57]^x[55]^x[47]^x[45]^x[36]^x[35]^x[34]^x[33];
	x_new[236]=x[376]^x[374]^x[370]^x[368]^x[366]^x[364]^x[359]^x[357]^x[355]^x[343]^x[337]^x[332]^x[331]^x[326]^x[320]^x[281]^x[280]^x[279]^x[275]^x[274]^x[273]^x[270]^x[268]^x[264]^x[263]^x[262]^x[237]^x[236]^x[226]^x[210]^x[208]^x[199]^x[197]^x[183]^x[172]^x[171]^x[160]^x[121]^x[120]^x[119]^x[110]^x[56]^x[54]^x[46]^x[44]^x[35]^x[34]^x[33]^x[32];
	x_new[235]=x[375]^x[374]^x[369]^x[368]^x[365]^x[358]^x[357]^x[354]^x[342]^x[336]^x[331]^x[325]^x[280]^x[279]^x[278]^x[274]^x[273]^x[272]^x[269]^x[267]^x[263]^x[262]^x[261]^x[236]^x[235]^x[225]^x[209]^x[208]^x[198]^x[197]^x[182]^x[171]^x[120]^x[119]^x[118]^x[109]^x[55]^x[54]^x[45]^x[34]^x[33]^x[32];
	x_new[234]=x[374]^x[368]^x[364]^x[362]^x[357]^x[353]^x[341]^x[335]^x[330]^x[324]^x[279]^x[278]^x[277]^x[273]^x[272]^x[271]^x[268]^x[266]^x[262]^x[261]^x[260]^x[235]^x[234]^x[224]^x[208]^x[197]^x[181]^x[170]^x[119]^x[118]^x[117]^x[108]^x[54]^x[44]^x[42]^x[33]^x[32];
	x_new[233]=x[381]^x[373]^x[372]^x[371]^x[363]^x[359]^x[352]^x[340]^x[334]^x[329]^x[323]^x[282]^x[278]^x[277]^x[276]^x[272]^x[271]^x[270]^x[267]^x[265]^x[261]^x[259]^x[255]^x[233]^x[180]^x[169]^x[118]^x[117]^x[116]^x[107]^x[53]^x[52]^x[51]^x[43]^x[41]^x[32];
	x_new[232]=x[383]^x[380]^x[372]^x[371]^x[370]^x[358]^x[339]^x[333]^x[328]^x[322]^x[277]^x[276]^x[275]^x[271]^x[270]^x[269]^x[266]^x[264]^x[260]^x[258]^x[254]^x[232]^x[179]^x[168]^x[117]^x[116]^x[115]^x[106]^x[63]^x[52]^x[50]^x[40];
	x_new[231]=x[382]^x[379]^x[371]^x[370]^x[369]^x[357]^x[338]^x[332]^x[327]^x[321]^x[276]^x[275]^x[274]^x[270]^x[269]^x[268]^x[265]^x[263]^x[259]^x[257]^x[253]^x[231]^x[178]^x[167]^x[138]^x[116]^x[115]^x[114]^x[105]^x[62]^x[51]^x[49]^x[39];
	x_new[230]=x[381]^x[378]^x[370]^x[369]^x[368]^x[356]^x[337]^x[331]^x[326]^x[320]^x[275]^x[274]^x[273]^x[269]^x[268]^x[267]^x[264]^x[262]^x[258]^x[256]^x[252]^x[230]^x[177]^x[166]^x[137]^x[115]^x[114]^x[113]^x[104]^x[61]^x[50]^x[48]^x[38];
	x_new[229]=x[380]^x[377]^x[374]^x[369]^x[367]^x[357]^x[355]^x[352]^x[336]^x[325]^x[278]^x[274]^x[273]^x[272]^x[263]^x[261]^x[256]^x[251]^x[229]^x[214]^x[192]^x[176]^x[165]^x[136]^x[114]^x[113]^x[112]^x[103]^x[60]^x[49]^x[47]^x[10];
	x_new[228]=x[379]^x[376]^x[373]^x[368]^x[366]^x[362]^x[356]^x[354]^x[335]^x[324]^x[273]^x[272]^x[271]^x[262]^x[260]^x[250]^x[228]^x[213]^x[202]^x[175]^x[164]^x[135]^x[113]^x[112]^x[111]^x[102]^x[59]^x[48]^x[46]^x[36]^x[9];
	x_new[227]=x[378]^x[375]^x[372]^x[367]^x[365]^x[361]^x[355]^x[353]^x[334]^x[323]^x[272]^x[271]^x[270]^x[261]^x[259]^x[249]^x[227]^x[212]^x[201]^x[174]^x[163]^x[134]^x[112]^x[111]^x[110]^x[101]^x[58]^x[47]^x[45]^x[35]^x[8];
	x_new[226]=x[377]^x[374]^x[371]^x[366]^x[364]^x[360]^x[354]^x[352]^x[333]^x[322]^x[271]^x[270]^x[269]^x[260]^x[258]^x[248]^x[226]^x[211]^x[200]^x[173]^x[162]^x[133]^x[111]^x[110]^x[109]^x[100]^x[57]^x[46]^x[44]^x[34]^x[7];
	x_new[225]=x[376]^x[370]^x[365]^x[363]^x[359]^x[353]^x[332]^x[321]^x[270]^x[269]^x[268]^x[259]^x[257]^x[247]^x[225]^x[210]^x[199]^x[172]^x[161]^x[110]^x[109]^x[108]^x[99]^x[56]^x[45]^x[43]^x[33]^x[6];
	x_new[224]=x[375]^x[369]^x[364]^x[363]^x[358]^x[331]^x[320]^x[269]^x[268]^x[267]^x[258]^x[256]^x[246]^x[224]^x[209]^x[198]^x[171]^x[160]^x[109]^x[108]^x[107]^x[98]^x[55]^x[44]^x[43]^x[5];
	x_new[223]=x[346]^x[345]^x[341]^x[336]^x[334]^x[332]^x[331]^x[330]^x[327]^x[325]^x[321]^x[319]^x[318]^x[313]^x[312]^x[309]^x[307]^x[303]^x[301]^x[298]^x[292]^x[284]^x[273]^x[255]^x[251]^x[250]^x[249]^x[247]^x[246]^x[245]^x[241]^x[239]^x[235]^x[234]^x[230]^x[229]^x[228]^x[225]^x[223]^x[213]^x[203]^x[192]^x[186]^x[185]^x[176]^x[174]^x[165]^x[159]^x[158]^x[149]^x[147]^x[138]^x[98]^x[87]^x[86]^x[85]^x[75]^x[74]^x[71]^x[65]^x[49]^x[43]^x[21]^x[20]^x[19]^x[12]^x[11]^x[1]^x[0];
	x_new[222]=x[350]^x[349]^x[338]^x[331]^x[330]^x[326]^x[320]^x[318]^x[317]^x[312]^x[311]^x[308]^x[306]^x[302]^x[300]^x[297]^x[291]^x[283]^x[272]^x[254]^x[248]^x[246]^x[245]^x[244]^x[240]^x[239]^x[238]^x[234]^x[233]^x[229]^x[228]^x[227]^x[224]^x[223]^x[222]^x[212]^x[158]^x[157]^x[148]^x[146]^x[137]^x[86]^x[85]^x[84]^x[74]^x[73]^x[70]^x[64]^x[48]^x[42]^x[30]^x[18]^x[11]^x[10]^x[0];
	x_new[221]=x[351]^x[349]^x[348]^x[337]^x[329]^x[325]^x[317]^x[316]^x[311]^x[310]^x[307]^x[305]^x[301]^x[299]^x[296]^x[290]^x[282]^x[271]^x[255]^x[253]^x[249]^x[247]^x[245]^x[244]^x[243]^x[239]^x[238]^x[237]^x[234]^x[233]^x[232]^x[228]^x[227]^x[226]^x[222]^x[221]^x[211]^x[157]^x[156]^x[147]^x[145]^x[136]^x[107]^x[96]^x[95]^x[85]^x[84]^x[83]^x[74]^x[73]^x[72]^x[69]^x[47]^x[41]^x[31]^x[29]^x[19]^x[17]^x[9];
	x_new[220]=x[350]^x[348]^x[347]^x[336]^x[328]^x[324]^x[316]^x[315]^x[310]^x[309]^x[306]^x[304]^x[300]^x[298]^x[295]^x[289]^x[281]^x[270]^x[254]^x[252]^x[248]^x[246]^x[244]^x[243]^x[242]^x[238]^x[237]^x[236]^x[233]^x[232]^x[231]^x[227]^x[226]^x[225]^x[221]^x[220]^x[210]^x[156]^x[155]^x[146]^x[144]^x[135]^x[106]^x[94]^x[84]^x[83]^x[82]^x[73]^x[72]^x[71]^x[68]^x[46]^x[40]^x[30]^x[28]^x[18]^x[16]^x[8];
	x_new[219]=x[349]^x[347]^x[346]^x[335]^x[327]^x[323]^x[315]^x[314]^x[309]^x[308]^x[305]^x[303]^x[299]^x[297]^x[294]^x[288]^x[280]^x[269]^x[253]^x[251]^x[247]^x[245]^x[243]^x[242]^x[241]^x[237]^x[236]^x[235]^x[232]^x[231]^x[230]^x[226]^x[225]^x[224]^x[220]^x[219]^x[209]^x[155]^x[154]^x[145]^x[143]^x[134]^x[105]^x[93]^x[83]^x[82]^x[81]^x[72]^x[71]^x[70]^x[67]^x[45]^x[39]^x[29]^x[27]^x[17]^x[15]^x[7];
	x_new[218]=x[383]^x[351]^x[350]^x[348]^x[344]^x[341]^x[340]^x[339]^x[335]^x[333]^x[331]^x[326]^x[322]^x[320]^x[319]^x[314]^x[313]^x[308]^x[307]^x[304]^x[302]^x[296]^x[293]^x[279]^x[268]^x[255]^x[252]^x[250]^x[245]^x[244]^x[242]^x[241]^x[240]^x[236]^x[231]^x[230]^x[229]^x[225]^x[224]^x[219]^x[218]^x[208]^x[191]^x[190]^x[181]^x[180]^x[179]^x[171]^x[160]^x[159]^x[154]^x[144]^x[142]^x[138]^x[133]^x[132]^x[125]^x[92]^x[82]^x[81]^x[80]^x[71]^x[70]^x[69]^x[66]^x[44]^x[38]^x[28]^x[16]^x[14]^x[6]^x[5];
	x_new[217]=x[382]^x[349]^x[347]^x[345]^x[344]^x[343]^x[340]^x[338]^x[334]^x[333]^x[332]^x[325]^x[321]^x[318]^x[313]^x[312]^x[307]^x[306]^x[303]^x[301]^x[295]^x[292]^x[278]^x[267]^x[255]^x[254]^x[251]^x[249]^x[245]^x[244]^x[243]^x[241]^x[240]^x[239]^x[235]^x[230]^x[229]^x[228]^x[224]^x[218]^x[217]^x[207]^x[189]^x[180]^x[178]^x[158]^x[153]^x[143]^x[141]^x[137]^x[132]^x[131]^x[124]^x[103]^x[91]^x[81]^x[80]^x[79]^x[70]^x[69]^x[68]^x[65]^x[43]^x[37]^x[27]^x[25]^x[15]^x[13]^x[5];
	x_new[216]=x[381]^x[348]^x[346]^x[344]^x[343]^x[342]^x[339]^x[337]^x[333]^x[332]^x[331]^x[324]^x[320]^x[317]^x[312]^x[311]^x[306]^x[305]^x[302]^x[300]^x[294]^x[291]^x[277]^x[266]^x[255]^x[254]^x[253]^x[250]^x[248]^x[244]^x[243]^x[242]^x[240]^x[239]^x[238]^x[229]^x[228]^x[227]^x[217]^x[216]^x[206]^x[188]^x[179]^x[177]^x[157]^x[152]^x[142]^x[140]^x[136]^x[131]^x[130]^x[123]^x[102]^x[90]^x[80]^x[79]^x[78]^x[69]^x[68]^x[67]^x[64]^x[42]^x[36]^x[26]^x[24]^x[14]^x[12]^x[4];
	x_new[215]=x[380]^x[347]^x[345]^x[343]^x[341]^x[338]^x[336]^x[332]^x[330]^x[323]^x[316]^x[311]^x[310]^x[305]^x[304]^x[301]^x[299]^x[293]^x[290]^x[276]^x[265]^x[254]^x[253]^x[252]^x[249]^x[247]^x[243]^x[242]^x[241]^x[239]^x[238]^x[237]^x[228]^x[227]^x[226]^x[216]^x[215]^x[205]^x[187]^x[178]^x[176]^x[156]^x[151]^x[141]^x[139]^x[135]^x[130]^x[129]^x[122]^x[89]^x[79]^x[78]^x[77]^x[68]^x[67]^x[66]^x[41]^x[35]^x[25]^x[23]^x[13]^x[11]^x[3];
	x_new[214]=x[379]^x[346]^x[344]^x[342]^x[340]^x[337]^x[335]^x[331]^x[329]^x[322]^x[315]^x[310]^x[309]^x[304]^x[303]^x[300]^x[298]^x[292]^x[289]^x[275]^x[264]^x[253]^x[252]^x[251]^x[248]^x[246]^x[242]^x[241]^x[240]^x[238]^x[237]^x[236]^x[227]^x[226]^x[225]^x[215]^x[214]^x[204]^x[186]^x[177]^x[175]^x[155]^x[150]^x[140]^x[138]^x[134]^x[129]^x[128]^x[121]^x[88]^x[78]^x[77]^x[76]^x[67]^x[66]^x[65]^x[40]^x[34]^x[24]^x[22]^x[12]^x[10]^x[2];
	x_new[213]=x[378]^x[345]^x[343]^x[341]^x[339]^x[336]^x[334]^x[331]^x[328]^x[321]^x[320]^x[314]^x[309]^x[308]^x[303]^x[302]^x[299]^x[297]^x[291]^x[288]^x[274]^x[263]^x[252]^x[251]^x[250]^x[247]^x[245]^x[241]^x[240]^x[239]^x[237]^x[236]^x[235]^x[226]^x[225]^x[224]^x[214]^x[213]^x[203]^x[185]^x[176]^x[174]^x[154]^x[149]^x[139]^x[137]^x[133]^x[128]^x[120]^x[87]^x[77]^x[76]^x[75]^x[66]^x[65]^x[64]^x[39]^x[33]^x[23]^x[21]^x[10]^x[9]^x[1]^x[0];
	x_new[212]=x[351]^x[350]^x[346]^x[345]^x[342]^x[340]^x[338]^x[334]^x[329]^x[320]^x[319]^x[313]^x[308]^x[307]^x[302]^x[301]^x[296]^x[290]^x[273]^x[262]^x[255]^x[251]^x[250]^x[249]^x[246]^x[244]^x[238]^x[236]^x[235]^x[229]^x[225]^x[224]^x[213]^x[212]^x[202]^x[186]^x[185]^x[174]^x[159]^x[148]^x[147]^x[136]^x[98]^x[95]^x[86]^x[76]^x[75]^x[65]^x[64]^x[38]^x[32]^x[31]^x[30]^x[22]^x[10]^x[9]^x[8]^x[0];
	x_new[211]=x[351]^x[349]^x[341]^x[338]^x[337]^x[330]^x[328]^x[327]^x[318]^x[312]^x[307]^x[306]^x[301]^x[300]^x[295]^x[289]^x[272]^x[261]^x[255]^x[254]^x[250]^x[249]^x[248]^x[245]^x[243]^x[239]^x[237]^x[235]^x[224]^x[212]^x[211]^x[201]^x[158]^x[147]^x[146]^x[135]^x[95]^x[94]^x[85]^x[75]^x[64]^x[37]^x[31]^x[29]^x[21]^x[19]^x[10]^x[9]^x[8]^x[7];
	x_new[210]=x[350]^x[348]^x[340]^x[337]^x[336]^x[329]^x[327]^x[326]^x[317]^x[311]^x[306]^x[305]^x[300]^x[299]^x[294]^x[288]^x[271]^x[260]^x[255]^x[254]^x[253]^x[249]^x[248]^x[247]^x[244]^x[242]^x[238]^x[236]^x[211]^x[210]^x[200]^x[157]^x[146]^x[145]^x[134]^x[95]^x[94]^x[93]^x[84]^x[36]^x[30]^x[28]^x[20]^x[18]^x[9]^x[8]^x[7]^x[6];
	x_new[209]=x[349]^x[347]^x[342]^x[341]^x[339]^x[330]^x[328]^x[326]^x[324]^x[320]^x[316]^x[310]^x[305]^x[304]^x[299]^x[293]^x[270]^x[259]^x[254]^x[253]^x[252]^x[248]^x[247]^x[246]^x[243]^x[241]^x[237]^x[235]^x[210]^x[209]^x[199]^x[182]^x[181]^x[170]^x[160]^x[156]^x[145]^x[144]^x[133]^x[94]^x[93]^x[92]^x[83]^x[35]^x[29]^x[27]^x[19]^x[17]^x[8]^x[7]^x[6]^x[5];
	x_new[208]=x[348]^x[346]^x[340]^x[338]^x[335]^x[329]^x[327]^x[325]^x[324]^x[323]^x[315]^x[309]^x[304]^x[303]^x[298]^x[292]^x[269]^x[258]^x[253]^x[252]^x[251]^x[247]^x[246]^x[245]^x[242]^x[240]^x[236]^x[234]^x[209]^x[208]^x[198]^x[180]^x[169]^x[155]^x[144]^x[143]^x[132]^x[93]^x[92]^x[91]^x[82]^x[34]^x[28]^x[26]^x[18]^x[16]^x[7]^x[6]^x[5]^x[4];
	x_new[207]=x[347]^x[345]^x[341]^x[339]^x[337]^x[335]^x[334]^x[330]^x[328]^x[326]^x[323]^x[322]^x[314]^x[308]^x[303]^x[302]^x[297]^x[291]^x[268]^x[257]^x[252]^x[251]^x[250]^x[246]^x[245]^x[244]^x[241]^x[239]^x[234]^x[233]^x[224]^x[208]^x[207]^x[197]^x[181]^x[179]^x[170]^x[168]^x[154]^x[143]^x[142]^x[131]^x[92]^x[91]^x[90]^x[81]^x[33]^x[27]^x[25]^x[17]^x[15]^x[6]^x[5]^x[4]^x[3];
	x_new[206]=x[346]^x[344]^x[340]^x[338]^x[336]^x[334]^x[333]^x[329]^x[327]^x[325]^x[322]^x[321]^x[313]^x[307]^x[302]^x[301]^x[296]^x[290]^x[267]^x[256]^x[251]^x[250]^x[249]^x[245]^x[244]^x[243]^x[240]^x[238]^x[234]^x[233]^x[232]^x[207]^x[206]^x[196]^x[180]^x[178]^x[169]^x[167]^x[153]^x[142]^x[141]^x[130]^x[91]^x[90]^x[89]^x[80]^x[32]^x[26]^x[24]^x[16]^x[14]^x[5]^x[4]^x[3]^x[2];
	x_new[205]=x[345]^x[343]^x[339]^x[337]^x[335]^x[333]^x[332]^x[328]^x[326]^x[324]^x[321]^x[320]^x[312]^x[306]^x[301]^x[300]^x[295]^x[289]^x[250]^x[249]^x[248]^x[244]^x[243]^x[242]^x[239]^x[237]^x[233]^x[232]^x[231]^x[206]^x[205]^x[195]^x[179]^x[177]^x[168]^x[166]^x[152]^x[141]^x[140]^x[129]^x[90]^x[89]^x[88]^x[79]^x[25]^x[23]^x[15]^x[13]^x[4]^x[3]^x[2]^x[1];
	x_new[204]=x[344]^x[342]^x[338]^x[336]^x[334]^x[332]^x[327]^x[325]^x[323]^x[311]^x[305]^x[300]^x[299]^x[294]^x[288]^x[249]^x[248]^x[247]^x[243]^x[242]^x[241]^x[238]^x[236]^x[232]^x[231]^x[230]^x[205]^x[204]^x[194]^x[178]^x[176]^x[167]^x[165]^x[151]^x[140]^x[139]^x[128]^x[89]^x[88]^x[87]^x[78]^x[24]^x[22]^x[14]^x[12]^x[3]^x[2]^x[1]^x[0];
	x_new[203]=x[343]^x[342]^x[337]^x[336]^x[333]^x[326]^x[325]^x[322]^x[310]^x[304]^x[299]^x[293]^x[248]^x[247]^x[246]^x[242]^x[241]^x[240]^x[237]^x[235]^x[231]^x[230]^x[229]^x[204]^x[203]^x[193]^x[177]^x[176]^x[166]^x[165]^x[150]^x[139]^x[88]^x[87]^x[86]^x[77]^x[23]^x[22]^x[13]^x[2]^x[1]^x[0];
	x_new[202]=x[342]^x[336]^x[332]^x[330]^x[325]^x[321]^x[309]^x[303]^x[298]^x[292]^x[247]^x[246]^x[245]^x[241]^x[240]^x[239]^x[236]^x[234]^x[230]^x[229]^x[228]^x[203]^x[202]^x[192]^x[176]^x[165]^x[149]^x[138]^x[87]^x[86]^x[85]^x[76]^x[22]^x[12]^x[10]^x[1]^x[0];
	x_new[201]=x[349]^x[341]^x[340]^x[339]^x[331]^x[327]^x[320]^x[308]^x[302]^x[297]^x[291]^x[250]^x[246]^x[245]^x[244]^x[240]^x[239]^x[238]^x[235]^x[233]^x[229]^x[227]^x[223]^x[201]^x[148]^x[137]^x[86]^x[85]^x[84]^x[75]^x[21]^x[20]^x[19]^x[11]^x[9]^x[0];
	x_new[200]=x[351]^x[348]^x[340]^x[339]^x[338]^x[326]^x[307]^x[301]^x[296]^x[290]^x[245]^x[244]^x[243]^x[239]^x[238]^x[237]^x[234]^x[232]^x[228]^x[226]^x[222]^x[200]^x[147]^x[136]^x[85]^x[84]^x[83]^x[74]^x[31]^x[20]^x[18]^x[8];
	x_new[199]=x[350]^x[347]^x[339]^x[338]^x[337]^x[325]^x[306]^x[300]^x[295]^x[289]^x[244]^x[243]^x[242]^x[238]^x[237]^x[236]^x[233]^x[231]^x[227]^x[225]^x[221]^x[199]^x[146]^x[135]^x[106]^x[84]^x[83]^x[82]^x[73]^x[30]^x[19]^x[17]^x[7];
	x_new[198]=x[349]^x[346]^x[338]^x[337]^x[336]^x[324]^x[305]^x[299]^x[294]^x[288]^x[243]^x[242]^x[241]^x[237]^x[236]^x[235]^x[232]^x[230]^x[226]^x[224]^x[220]^x[198]^x[145]^x[134]^x[105]^x[83]^x[82]^x[81]^x[72]^x[29]^x[18]^x[16]^x[6];
	x_new[197]=x[373]^x[362]^x[348]^x[345]^x[342]^x[337]^x[335]^x[325]^x[323]^x[320]^x[304]^x[293]^x[246]^x[242]^x[241]^x[240]^x[231]^x[229]^x[224]^x[219]^x[197]^x[182]^x[160]^x[144]^x[138]^x[133]^x[132]^x[104]^x[82]^x[81]^x[80]^x[71]^x[28]^x[17]^x[15];
	x_new[196]=x[372]^x[361]^x[347]^x[344]^x[341]^x[336]^x[334]^x[330]^x[324]^x[322]^x[303]^x[292]^x[241]^x[240]^x[239]^x[230]^x[228]^x[218]^x[196]^x[181]^x[170]^x[143]^x[137]^x[132]^x[131]^x[103]^x[81]^x[80]^x[79]^x[70]^x[27]^x[16]^x[14]^x[4];
	x_new[195]=x[371]^x[360]^x[346]^x[343]^x[340]^x[335]^x[333]^x[329]^x[323]^x[321]^x[302]^x[291]^x[240]^x[239]^x[238]^x[229]^x[227]^x[217]^x[195]^x[180]^x[169]^x[142]^x[136]^x[131]^x[130]^x[102]^x[80]^x[79]^x[78]^x[69]^x[26]^x[15]^x[13]^x[3];
	x_new[194]=x[370]^x[359]^x[345]^x[342]^x[339]^x[334]^x[332]^x[328]^x[322]^x[320]^x[301]^x[290]^x[239]^x[238]^x[237]^x[228]^x[226]^x[216]^x[194]^x[179]^x[168]^x[141]^x[135]^x[130]^x[129]^x[101]^x[79]^x[78]^x[77]^x[68]^x[25]^x[14]^x[12]^x[2];
	x_new[193]=x[369]^x[358]^x[344]^x[338]^x[333]^x[331]^x[327]^x[321]^x[300]^x[289]^x[238]^x[237]^x[236]^x[227]^x[225]^x[215]^x[193]^x[178]^x[167]^x[140]^x[134]^x[129]^x[128]^x[78]^x[77]^x[76]^x[67]^x[24]^x[13]^x[11]^x[1];
	x_new[192]=x[368]^x[357]^x[343]^x[337]^x[332]^x[331]^x[326]^x[299]^x[288]^x[237]^x[236]^x[235]^x[226]^x[224]^x[214]^x[192]^x[177]^x[166]^x[139]^x[133]^x[128]^x[77]^x[76]^x[75]^x[66]^x[23]^x[12]^x[11];
	x_new[191]=x[383]^x[382]^x[375]^x[374]^x[373]^x[372]^x[371]^x[363]^x[353]^x[314]^x[313]^x[309]^x[304]^x[302]^x[300]^x[299]^x[298]^x[295]^x[293]^x[289]^x[287]^x[286]^x[281]^x[280]^x[277]^x[275]^x[271]^x[269]^x[266]^x[260]^x[252]^x[241]^x[223]^x[219]^x[218]^x[217]^x[215]^x[214]^x[213]^x[209]^x[207]^x[203]^x[202]^x[198]^x[197]^x[196]^x[193]^x[191]^x[181]^x[171]^x[160]^x[154]^x[153]^x[149]^x[148]^x[147]^x[144]^x[143]^x[141]^x[140]^x[139]^x[134]^x[129]^x[128]^x[127]^x[126]^x[117]^x[115]^x[106]^x[66]^x[55]^x[54]^x[53]^x[43]^x[42]^x[39]^x[33]^x[17]^x[11];
	x_new[190]=x[382]^x[381]^x[374]^x[373]^x[372]^x[370]^x[362]^x[361]^x[352]^x[318]^x[317]^x[306]^x[299]^x[298]^x[294]^x[288]^x[286]^x[285]^x[280]^x[279]^x[276]^x[274]^x[270]^x[268]^x[265]^x[259]^x[251]^x[240]^x[222]^x[216]^x[214]^x[213]^x[212]^x[208]^x[207]^x[206]^x[202]^x[201]^x[197]^x[196]^x[195]^x[192]^x[191]^x[190]^x[180]^x[158]^x[152]^x[146]^x[140]^x[139]^x[138]^x[133]^x[132]^x[128]^x[126]^x[125]^x[116]^x[114]^x[105]^x[54]^x[53]^x[52]^x[42]^x[41]^x[38]^x[32]^x[16]^x[10];
	x_new[189]=x[383]^x[382]^x[381]^x[380]^x[373]^x[372]^x[369]^x[362]^x[361]^x[360]^x[319]^x[317]^x[316]^x[305]^x[297]^x[293]^x[285]^x[284]^x[279]^x[278]^x[275]^x[273]^x[269]^x[267]^x[264]^x[258]^x[250]^x[239]^x[223]^x[221]^x[217]^x[215]^x[213]^x[212]^x[211]^x[207]^x[206]^x[205]^x[202]^x[201]^x[200]^x[196]^x[195]^x[194]^x[190]^x[189]^x[179]^x[159]^x[157]^x[153]^x[151]^x[147]^x[145]^x[141]^x[139]^x[137]^x[131]^x[125]^x[124]^x[115]^x[113]^x[104]^x[75]^x[64]^x[63]^x[53]^x[52]^x[51]^x[42]^x[41]^x[40]^x[37]^x[15]^x[9];
	x_new[188]=x[382]^x[381]^x[380]^x[379]^x[372]^x[371]^x[368]^x[361]^x[360]^x[359]^x[318]^x[316]^x[315]^x[304]^x[296]^x[292]^x[284]^x[283]^x[278]^x[277]^x[274]^x[272]^x[268]^x[266]^x[263]^x[257]^x[249]^x[238]^x[222]^x[220]^x[216]^x[214]^x[212]^x[211]^x[210]^x[206]^x[205]^x[204]^x[201]^x[200]^x[199]^x[195]^x[194]^x[193]^x[189]^x[188]^x[178]^x[158]^x[156]^x[152]^x[150]^x[146]^x[144]^x[140]^x[138]^x[136]^x[130]^x[124]^x[123]^x[114]^x[112]^x[103]^x[74]^x[62]^x[52]^x[51]^x[50]^x[41]^x[40]^x[39]^x[36]^x[14]^x[8];
	x_new[187]=x[381]^x[380]^x[379]^x[378]^x[371]^x[370]^x[367]^x[360]^x[359]^x[358]^x[317]^x[315]^x[314]^x[303]^x[295]^x[291]^x[283]^x[282]^x[277]^x[276]^x[273]^x[271]^x[267]^x[265]^x[262]^x[256]^x[248]^x[237]^x[221]^x[219]^x[215]^x[213]^x[211]^x[210]^x[209]^x[205]^x[204]^x[203]^x[200]^x[199]^x[198]^x[194]^x[193]^x[192]^x[188]^x[187]^x[177]^x[157]^x[155]^x[151]^x[149]^x[145]^x[143]^x[139]^x[137]^x[135]^x[129]^x[123]^x[122]^x[113]^x[111]^x[102]^x[73]^x[61]^x[51]^x[50]^x[49]^x[40]^x[39]^x[38]^x[35]^x[13]^x[7];
	x_new[186]=x[380]^x[379]^x[377]^x[370]^x[369]^x[366]^x[359]^x[358]^x[357]^x[351]^x[319]^x[318]^x[316]^x[312]^x[309]^x[308]^x[307]^x[303]^x[301]^x[299]^x[294]^x[290]^x[288]^x[287]^x[282]^x[281]^x[276]^x[275]^x[272]^x[270]^x[264]^x[261]^x[247]^x[236]^x[223]^x[220]^x[218]^x[213]^x[212]^x[210]^x[209]^x[208]^x[204]^x[199]^x[198]^x[197]^x[193]^x[192]^x[187]^x[186]^x[176]^x[159]^x[158]^x[156]^x[150]^x[149]^x[148]^x[147]^x[144]^x[142]^x[139]^x[138]^x[136]^x[134]^x[133]^x[127]^x[122]^x[112]^x[110]^x[106]^x[101]^x[100]^x[93]^x[60]^x[50]^x[49]^x[48]^x[39]^x[38]^x[37]^x[34]^x[12]^x[6];
	x_new[185]=x[379]^x[378]^x[377]^x[376]^x[369]^x[368]^x[365]^x[358]^x[357]^x[356]^x[350]^x[317]^x[315]^x[313]^x[312]^x[311]^x[308]^x[306]^x[302]^x[301]^x[300]^x[293]^x[289]^x[286]^x[281]^x[280]^x[275]^x[274]^x[271]^x[269]^x[263]^x[260]^x[246]^x[235]^x[223]^x[222]^x[219]^x[217]^x[213]^x[212]^x[211]^x[209]^x[208]^x[207]^x[203]^x[198]^x[197]^x[196]^x[192]^x[186]^x[185]^x[175]^x[157]^x[155]^x[153]^x[149]^x[148]^x[147]^x[146]^x[143]^x[141]^x[137]^x[135]^x[133]^x[126]^x[121]^x[111]^x[109]^x[105]^x[100]^x[99]^x[92]^x[71]^x[59]^x[49]^x[48]^x[47]^x[38]^x[37]^x[36]^x[33]^x[11]^x[5];
	x_new[184]=x[378]^x[377]^x[376]^x[375]^x[368]^x[367]^x[364]^x[357]^x[356]^x[355]^x[349]^x[316]^x[314]^x[312]^x[311]^x[310]^x[307]^x[305]^x[301]^x[300]^x[299]^x[292]^x[288]^x[285]^x[280]^x[279]^x[274]^x[273]^x[270]^x[268]^x[262]^x[259]^x[245]^x[234]^x[223]^x[222]^x[221]^x[218]^x[216]^x[212]^x[211]^x[210]^x[208]^x[207]^x[206]^x[197]^x[196]^x[195]^x[185]^x[184]^x[174]^x[156]^x[154]^x[152]^x[148]^x[147]^x[146]^x[145]^x[142]^x[140]^x[136]^x[134]^x[132]^x[125]^x[120]^x[110]^x[108]^x[104]^x[99]^x[98]^x[91]^x[70]^x[58]^x[48]^x[47]^x[46]^x[37]^x[36]^x[35]^x[32]^x[10]^x[4];
	x_new[183]=x[377]^x[376]^x[375]^x[374]^x[367]^x[366]^x[363]^x[356]^x[355]^x[354]^x[348]^x[315]^x[313]^x[311]^x[309]^x[306]^x[304]^x[300]^x[298]^x[291]^x[284]^x[279]^x[278]^x[273]^x[272]^x[269]^x[267]^x[261]^x[258]^x[244]^x[233]^x[222]^x[221]^x[220]^x[217]^x[215]^x[211]^x[210]^x[209]^x[207]^x[206]^x[205]^x[196]^x[195]^x[194]^x[184]^x[183]^x[173]^x[155]^x[153]^x[151]^x[147]^x[146]^x[145]^x[144]^x[141]^x[139]^x[135]^x[133]^x[131]^x[124]^x[119]^x[109]^x[107]^x[103]^x[98]^x[97]^x[90]^x[57]^x[47]^x[46]^x[45]^x[36]^x[35]^x[34]^x[9]^x[3];
	x_new[182]=x[376]^x[375]^x[374]^x[373]^x[366]^x[365]^x[362]^x[355]^x[354]^x[353]^x[347]^x[314]^x[312]^x[310]^x[308]^x[305]^x[303]^x[299]^x[297]^x[290]^x[283]^x[278]^x[277]^x[272]^x[271]^x[268]^x[266]^x[260]^x[257]^x[243]^x[232]^x[221]^x[220]^x[219]^x[216]^x[214]^x[210]^x[209]^x[208]^x[206]^x[205]^x[204]^x[195]^x[194]^x[193]^x[183]^x[182]^x[172]^x[154]^x[152]^x[150]^x[146]^x[145]^x[144]^x[143]^x[140]^x[138]^x[134]^x[132]^x[130]^x[123]^x[118]^x[108]^x[106]^x[102]^x[97]^x[96]^x[89]^x[56]^x[46]^x[45]^x[44]^x[35]^x[34]^x[33]^x[8]^x[2];
	x_new[181]=x[375]^x[372]^x[365]^x[364]^x[362]^x[361]^x[354]^x[353]^x[346]^x[313]^x[311]^x[309]^x[307]^x[304]^x[302]^x[299]^x[296]^x[289]^x[288]^x[282]^x[277]^x[276]^x[271]^x[270]^x[267]^x[265]^x[259]^x[256]^x[242]^x[231]^x[220]^x[219]^x[218]^x[215]^x[213]^x[209]^x[208]^x[207]^x[205]^x[204]^x[203]^x[194]^x[193]^x[192]^x[182]^x[181]^x[171]^x[153]^x[151]^x[149]^x[145]^x[144]^x[143]^x[142]^x[138]^x[137]^x[132]^x[131]^x[129]^x[128]^x[122]^x[117]^x[107]^x[105]^x[101]^x[96]^x[88]^x[55]^x[45]^x[44]^x[43]^x[34]^x[33]^x[32]^x[7]^x[1];
	x_new[180]=x[383]^x[382]^x[374]^x[371]^x[364]^x[363]^x[360]^x[353]^x[352]^x[319]^x[318]^x[314]^x[313]^x[310]^x[308]^x[306]^x[302]^x[297]^x[288]^x[287]^x[281]^x[276]^x[275]^x[270]^x[269]^x[264]^x[258]^x[241]^x[230]^x[223]^x[219]^x[218]^x[217]^x[214]^x[212]^x[206]^x[204]^x[203]^x[197]^x[193]^x[192]^x[181]^x[180]^x[170]^x[159]^x[158]^x[154]^x[152]^x[150]^x[144]^x[142]^x[138]^x[137]^x[136]^x[132]^x[131]^x[130]^x[128]^x[127]^x[116]^x[115]^x[104]^x[66]^x[63]^x[54]^x[44]^x[43]^x[33]^x[32]^x[6]^x[0];
	x_new[179]=x[383]^x[382]^x[381]^x[373]^x[372]^x[371]^x[370]^x[363]^x[361]^x[359]^x[352]^x[319]^x[317]^x[309]^x[306]^x[305]^x[298]^x[296]^x[295]^x[286]^x[280]^x[275]^x[274]^x[269]^x[268]^x[263]^x[257]^x[240]^x[229]^x[223]^x[222]^x[218]^x[217]^x[216]^x[213]^x[211]^x[207]^x[205]^x[203]^x[192]^x[180]^x[179]^x[169]^x[159]^x[157]^x[153]^x[151]^x[149]^x[147]^x[143]^x[141]^x[138]^x[137]^x[136]^x[135]^x[132]^x[131]^x[130]^x[129]^x[126]^x[115]^x[114]^x[103]^x[63]^x[62]^x[53]^x[43]^x[32]^x[5];
	x_new[178]=x[383]^x[382]^x[381]^x[380]^x[372]^x[371]^x[370]^x[369]^x[360]^x[358]^x[318]^x[316]^x[308]^x[305]^x[304]^x[297]^x[295]^x[294]^x[285]^x[279]^x[274]^x[273]^x[268]^x[267]^x[262]^x[256]^x[239]^x[228]^x[223]^x[222]^x[221]^x[217]^x[216]^x[215]^x[212]^x[210]^x[206]^x[204]^x[179]^x[178]^x[168]^x[158]^x[156]^x[152]^x[150]^x[148]^x[146]^x[142]^x[140]^x[137]^x[136]^x[135]^x[134]^x[131]^x[130]^x[129]^x[128]^x[125]^x[114]^x[113]^x[102]^x[63]^x[62]^x[61]^x[52]^x[4];
	x_new[177]=x[382]^x[381]^x[380]^x[379]^x[371]^x[370]^x[369]^x[368]^x[359]^x[357]^x[317]^x[315]^x[310]^x[309]^x[307]^x[298]^x[296]^x[294]^x[292]^x[288]^x[284]^x[278]^x[273]^x[272]^x[267]^x[261]^x[238]^x[227]^x[222]^x[221]^x[220]^x[216]^x[215]^x[214]^x[211]^x[209]^x[205]^x[203]^x[178]^x[177]^x[167]^x[157]^x[155]^x[151]^x[150]^x[147]^x[145]^x[141]^x[139]^x[138]^x[136]^x[135]^x[134]^x[133]^x[130]^x[129]^x[124]^x[113]^x[112]^x[101]^x[62]^x[61]^x[60]^x[51]^x[3];
	x_new[176]=x[381]^x[380]^x[379]^x[378]^x[370]^x[369]^x[368]^x[367]^x[358]^x[356]^x[316]^x[314]^x[308]^x[306]^x[303]^x[297]^x[295]^x[293]^x[292]^x[291]^x[283]^x[277]^x[272]^x[271]^x[266]^x[260]^x[237]^x[226]^x[221]^x[220]^x[219]^x[215]^x[214]^x[213]^x[210]^x[208]^x[204]^x[202]^x[177]^x[176]^x[166]^x[156]^x[154]^x[150]^x[146]^x[144]^x[140]^x[138]^x[137]^x[135]^x[134]^x[133]^x[132]^x[129]^x[128]^x[123]^x[112]^x[111]^x[100]^x[61]^x[60]^x[59]^x[50]^x[2];
	x_new[175]=x[380]^x[379]^x[378]^x[377]^x[369]^x[368]^x[367]^x[366]^x[357]^x[355]^x[315]^x[313]^x[309]^x[307]^x[305]^x[303]^x[302]^x[298]^x[296]^x[294]^x[291]^x[290]^x[282]^x[276]^x[271]^x[270]^x[265]^x[259]^x[236]^x[225]^x[220]^x[219]^x[218]^x[214]^x[213]^x[212]^x[209]^x[207]^x[202]^x[201]^x[192]^x[176]^x[175]^x[165]^x[155]^x[153]^x[145]^x[143]^x[139]^x[138]^x[137]^x[136]^x[134]^x[133]^x[132]^x[131]^x[128]^x[122]^x[111]^x[110]^x[99]^x[60]^x[59]^x[58]^x[49]^x[1];
	x_new[174]=x[379]^x[378]^x[377]^x[376]^x[368]^x[367]^x[366]^x[365]^x[356]^x[354]^x[314]^x[312]^x[308]^x[306]^x[304]^x[302]^x[301]^x[297]^x[295]^x[293]^x[290]^x[289]^x[281]^x[275]^x[270]^x[269]^x[264]^x[258]^x[235]^x[224]^x[219]^x[218]^x[217]^x[213]^x[212]^x[211]^x[208]^x[206]^x[202]^x[201]^x[200]^x[175]^x[174]^x[164]^x[154]^x[152]^x[144]^x[142]^x[138]^x[137]^x[136]^x[135]^x[133]^x[132]^x[131]^x[130]^x[121]^x[110]^x[109]^x[98]^x[59]^x[58]^x[57]^x[48]^x[0];
	x_new[173]=x[378]^x[377]^x[376]^x[375]^x[367]^x[366]^x[365]^x[364]^x[355]^x[353]^x[313]^x[311]^x[307]^x[305]^x[303]^x[301]^x[300]^x[296]^x[294]^x[292]^x[289]^x[288]^x[280]^x[274]^x[269]^x[268]^x[263]^x[257]^x[218]^x[217]^x[216]^x[212]^x[211]^x[210]^x[207]^x[205]^x[201]^x[200]^x[199]^x[174]^x[173]^x[163]^x[153]^x[151]^x[143]^x[141]^x[137]^x[136]^x[135]^x[134]^x[132]^x[131]^x[130]^x[129]^x[120]^x[109]^x[108]^x[97]^x[58]^x[57]^x[56]^x[47];
	x_new[172]=x[377]^x[376]^x[375]^x[374]^x[366]^x[365]^x[364]^x[363]^x[354]^x[352]^x[312]^x[310]^x[306]^x[304]^x[302]^x[300]^x[295]^x[293]^x[291]^x[279]^x[273]^x[268]^x[267]^x[262]^x[256]^x[217]^x[216]^x[215]^x[211]^x[210]^x[209]^x[206]^x[204]^x[200]^x[199]^x[198]^x[173]^x[172]^x[162]^x[152]^x[150]^x[142]^x[140]^x[136]^x[135]^x[134]^x[133]^x[131]^x[130]^x[129]^x[128]^x[119]^x[108]^x[107]^x[96]^x[57]^x[56]^x[55]^x[46];
	x_new[171]=x[376]^x[375]^x[374]^x[365]^x[363]^x[352]^x[311]^x[310]^x[305]^x[304]^x[301]^x[294]^x[293]^x[290]^x[278]^x[272]^x[267]^x[261]^x[216]^x[215]^x[214]^x[210]^x[209]^x[208]^x[205]^x[203]^x[199]^x[198]^x[197]^x[172]^x[171]^x[161]^x[151]^x[150]^x[141]^x[135]^x[134]^x[133]^x[130]^x[129]^x[128]^x[118]^x[107]^x[56]^x[55]^x[54]^x[45];
	x_new[170]=x[375]^x[374]^x[373]^x[364]^x[363]^x[362]^x[352]^x[310]^x[304]^x[300]^x[298]^x[293]^x[289]^x[277]^x[271]^x[266]^x[260]^x[215]^x[214]^x[213]^x[209]^x[208]^x[207]^x[204]^x[202]^x[198]^x[197]^x[196]^x[171]^x[170]^x[160]^x[150]^x[140]^x[138]^x[134]^x[133]^x[132]^x[129]^x[128]^x[117]^x[106]^x[55]^x[54]^x[53]^x[44];
	x_new[169]=x[383]^x[382]^x[374]^x[373]^x[371]^x[363]^x[361]^x[317]^x[309]^x[308]^x[307]^x[299]^x[295]^x[288]^x[276]^x[270]^x[265]^x[259]^x[218]^x[214]^x[213]^x[212]^x[208]^x[207]^x[206]^x[203]^x[201]^x[197]^x[195]^x[191]^x[169]^x[149]^x[148]^x[147]^x[143]^x[142]^x[141]^x[139]^x[137]^x[133]^x[131]^x[128]^x[116]^x[105]^x[54]^x[53]^x[52]^x[43];
	x_new[168]=x[381]^x[373]^x[372]^x[371]^x[370]^x[362]^x[360]^x[319]^x[316]^x[308]^x[307]^x[306]^x[294]^x[275]^x[269]^x[264]^x[258]^x[213]^x[212]^x[211]^x[207]^x[206]^x[205]^x[202]^x[200]^x[196]^x[194]^x[190]^x[168]^x[159]^x[153]^x[148]^x[146]^x[142]^x[140]^x[136]^x[130]^x[115]^x[104]^x[53]^x[52]^x[51]^x[42];
	x_new[167]=x[380]^x[372]^x[371]^x[370]^x[369]^x[361]^x[359]^x[318]^x[315]^x[307]^x[306]^x[305]^x[293]^x[274]^x[268]^x[263]^x[257]^x[212]^x[211]^x[210]^x[206]^x[205]^x[204]^x[201]^x[199]^x[195]^x[193]^x[189]^x[167]^x[158]^x[152]^x[147]^x[145]^x[141]^x[139]^x[135]^x[129]^x[114]^x[103]^x[74]^x[52]^x[51]^x[50]^x[41];
	x_new[166]=x[379]^x[371]^x[370]^x[369]^x[368]^x[360]^x[358]^x[317]^x[314]^x[306]^x[305]^x[304]^x[292]^x[273]^x[267]^x[262]^x[256]^x[211]^x[210]^x[209]^x[205]^x[204]^x[203]^x[200]^x[198]^x[194]^x[192]^x[188]^x[166]^x[157]^x[151]^x[146]^x[144]^x[140]^x[138]^x[134]^x[128]^x[113]^x[102]^x[73]^x[51]^x[50]^x[49]^x[40];
	x_new[165]=x[378]^x[370]^x[369]^x[367]^x[359]^x[341]^x[330]^x[316]^x[313]^x[310]^x[305]^x[303]^x[293]^x[291]^x[288]^x[272]^x[261]^x[214]^x[210]^x[209]^x[208]^x[199]^x[197]^x[192]^x[187]^x[165]^x[156]^x[145]^x[143]^x[139]^x[137]^x[128]^x[112]^x[106]^x[101]^x[100]^x[72]^x[50]^x[49]^x[48]^x[39];
	x_new[164]=x[377]^x[369]^x[368]^x[367]^x[366]^x[358]^x[356]^x[340]^x[329]^x[315]^x[312]^x[309]^x[304]^x[302]^x[298]^x[292]^x[290]^x[271]^x[260]^x[209]^x[208]^x[207]^x[198]^x[196]^x[186]^x[164]^x[155]^x[144]^x[142]^x[136]^x[132]^x[111]^x[105]^x[100]^x[99]^x[71]^x[49]^x[48]^x[47]^x[38];
	x_new[163]=x[376]^x[368]^x[367]^x[366]^x[365]^x[357]^x[355]^x[339]^x[328]^x[314]^x[311]^x[308]^x[303]^x[301]^x[297]^x[291]^x[289]^x[270]^x[259]^x[208]^x[207]^x[206]^x[197]^x[195]^x[185]^x[163]^x[154]^x[143]^x[141]^x[135]^x[131]^x[110]^x[104]^x[99]^x[98]^x[70]^x[48]^x[47]^x[46]^x[37];
	x_new[162]=x[375]^x[367]^x[366]^x[365]^x[364]^x[356]^x[354]^x[338]^x[327]^x[313]^x[310]^x[307]^x[302]^x[300]^x[296]^x[290]^x[288]^x[269]^x[258]^x[207]^x[206]^x[205]^x[196]^x[194]^x[184]^x[162]^x[153]^x[142]^x[140]^x[134]^x[130]^x[109]^x[103]^x[98]^x[97]^x[69]^x[47]^x[46]^x[45]^x[36];
	x_new[161]=x[374]^x[366]^x[365]^x[364]^x[363]^x[355]^x[353]^x[337]^x[326]^x[312]^x[306]^x[301]^x[299]^x[295]^x[289]^x[268]^x[257]^x[206]^x[205]^x[204]^x[195]^x[193]^x[183]^x[161]^x[152]^x[141]^x[139]^x[133]^x[129]^x[108]^x[102]^x[97]^x[96]^x[46]^x[45]^x[44]^x[35];
	x_new[160]=x[374]^x[365]^x[364]^x[363]^x[354]^x[336]^x[325]^x[311]^x[305]^x[300]^x[299]^x[294]^x[267]^x[256]^x[205]^x[204]^x[203]^x[194]^x[192]^x[182]^x[160]^x[151]^x[140]^x[139]^x[133]^x[107]^x[101]^x[96]^x[45]^x[44]^x[43]^x[34];
	x_new[159]=x[380]^x[374]^x[369]^x[363]^x[351]^x[350]^x[343]^x[342]^x[341]^x[340]^x[339]^x[331]^x[321]^x[282]^x[281]^x[277]^x[272]^x[270]^x[268]^x[267]^x[266]^x[263]^x[261]^x[257]^x[255]^x[254]^x[249]^x[248]^x[245]^x[243]^x[239]^x[237]^x[234]^x[228]^x[220]^x[209]^x[191]^x[187]^x[186]^x[185]^x[183]^x[182]^x[181]^x[177]^x[175]^x[171]^x[170]^x[166]^x[165]^x[164]^x[161]^x[159]^x[149]^x[145]^x[139]^x[133]^x[128]^x[122]^x[121]^x[117]^x[116]^x[115]^x[112]^x[111]^x[109]^x[108]^x[107]^x[102]^x[97]^x[96]^x[95]^x[94]^x[85]^x[83]^x[74]^x[34]^x[23]^x[22]^x[21]^x[11]^x[10]^x[7]^x[1];
	x_new[158]=x[379]^x[373]^x[368]^x[362]^x[350]^x[349]^x[342]^x[341]^x[340]^x[338]^x[330]^x[329]^x[320]^x[286]^x[285]^x[274]^x[267]^x[266]^x[262]^x[256]^x[254]^x[253]^x[248]^x[247]^x[244]^x[242]^x[238]^x[236]^x[233]^x[227]^x[219]^x[208]^x[190]^x[184]^x[182]^x[181]^x[180]^x[176]^x[175]^x[174]^x[170]^x[169]^x[165]^x[164]^x[163]^x[160]^x[159]^x[158]^x[148]^x[144]^x[132]^x[126]^x[120]^x[114]^x[108]^x[107]^x[106]^x[101]^x[100]^x[96]^x[94]^x[93]^x[84]^x[82]^x[73]^x[22]^x[21]^x[20]^x[10]^x[9]^x[6]^x[0];
	x_new[157]=x[378]^x[372]^x[367]^x[361]^x[351]^x[350]^x[349]^x[348]^x[341]^x[340]^x[337]^x[330]^x[329]^x[328]^x[287]^x[285]^x[284]^x[273]^x[265]^x[261]^x[253]^x[252]^x[247]^x[246]^x[243]^x[241]^x[237]^x[235]^x[232]^x[226]^x[218]^x[207]^x[191]^x[189]^x[185]^x[183]^x[181]^x[180]^x[179]^x[175]^x[174]^x[173]^x[170]^x[169]^x[168]^x[164]^x[163]^x[162]^x[158]^x[157]^x[147]^x[143]^x[131]^x[127]^x[125]^x[121]^x[119]^x[115]^x[113]^x[109]^x[107]^x[105]^x[99]^x[93]^x[92]^x[83]^x[81]^x[72]^x[43]^x[32]^x[31]^x[21]^x[20]^x[19]^x[10]^x[9]^x[8]^x[5];
	x_new[156]=x[377]^x[371]^x[366]^x[360]^x[350]^x[349]^x[348]^x[347]^x[340]^x[339]^x[336]^x[329]^x[328]^x[327]^x[286]^x[284]^x[283]^x[272]^x[264]^x[260]^x[252]^x[251]^x[246]^x[245]^x[242]^x[240]^x[236]^x[234]^x[231]^x[225]^x[217]^x[206]^x[190]^x[188]^x[184]^x[182]^x[180]^x[179]^x[178]^x[174]^x[173]^x[172]^x[169]^x[168]^x[167]^x[163]^x[162]^x[161]^x[157]^x[156]^x[146]^x[142]^x[130]^x[126]^x[124]^x[120]^x[118]^x[114]^x[112]^x[108]^x[106]^x[104]^x[98]^x[92]^x[91]^x[82]^x[80]^x[71]^x[42]^x[30]^x[20]^x[19]^x[18]^x[9]^x[8]^x[7]^x[4];
	x_new[155]=x[376]^x[370]^x[365]^x[359]^x[349]^x[348]^x[347]^x[346]^x[339]^x[338]^x[335]^x[328]^x[327]^x[326]^x[285]^x[283]^x[282]^x[271]^x[263]^x[259]^x[251]^x[250]^x[245]^x[244]^x[241]^x[239]^x[235]^x[233]^x[230]^x[224]^x[216]^x[205]^x[189]^x[187]^x[183]^x[181]^x[179]^x[178]^x[177]^x[173]^x[172]^x[171]^x[168]^x[167]^x[166]^x[162]^x[161]^x[160]^x[156]^x[155]^x[145]^x[141]^x[129]^x[125]^x[123]^x[119]^x[117]^x[113]^x[111]^x[107]^x[105]^x[103]^x[97]^x[91]^x[90]^x[81]^x[79]^x[70]^x[41]^x[29]^x[19]^x[18]^x[17]^x[8]^x[7]^x[6]^x[3];
	x_new[154]=x[375]^x[369]^x[364]^x[358]^x[348]^x[347]^x[345]^x[338]^x[337]^x[334]^x[327]^x[326]^x[325]^x[319]^x[287]^x[286]^x[284]^x[280]^x[277]^x[276]^x[275]^x[271]^x[269]^x[267]^x[262]^x[258]^x[256]^x[255]^x[250]^x[249]^x[244]^x[243]^x[240]^x[238]^x[232]^x[229]^x[215]^x[204]^x[191]^x[188]^x[186]^x[181]^x[180]^x[178]^x[177]^x[176]^x[172]^x[167]^x[166]^x[165]^x[161]^x[160]^x[155]^x[154]^x[144]^x[140]^x[128]^x[127]^x[126]^x[124]^x[118]^x[117]^x[116]^x[115]^x[112]^x[110]^x[107]^x[106]^x[104]^x[102]^x[101]^x[95]^x[90]^x[80]^x[78]^x[74]^x[69]^x[68]^x[61]^x[28]^x[18]^x[17]^x[16]^x[7]^x[6]^x[5]^x[2];
	x_new[153]=x[374]^x[368]^x[363]^x[357]^x[347]^x[346]^x[345]^x[344]^x[337]^x[336]^x[333]^x[326]^x[325]^x[324]^x[318]^x[285]^x[283]^x[281]^x[280]^x[279]^x[276]^x[274]^x[270]^x[269]^x[268]^x[261]^x[257]^x[254]^x[249]^x[248]^x[243]^x[242]^x[239]^x[237]^x[231]^x[228]^x[214]^x[203]^x[191]^x[190]^x[187]^x[185]^x[181]^x[180]^x[179]^x[177]^x[176]^x[175]^x[171]^x[166]^x[165]^x[164]^x[160]^x[154]^x[153]^x[143]^x[139]^x[125]^x[123]^x[121]^x[117]^x[116]^x[115]^x[114]^x[111]^x[109]^x[105]^x[103]^x[101]^x[94]^x[89]^x[79]^x[77]^x[73]^x[68]^x[67]^x[60]^x[39]^x[27]^x[17]^x[16]^x[15]^x[6]^x[5]^x[4]^x[1];
	x_new[152]=x[373]^x[367]^x[362]^x[356]^x[346]^x[345]^x[344]^x[343]^x[336]^x[335]^x[332]^x[325]^x[324]^x[323]^x[317]^x[284]^x[282]^x[280]^x[279]^x[278]^x[275]^x[273]^x[269]^x[268]^x[267]^x[260]^x[256]^x[253]^x[248]^x[247]^x[242]^x[241]^x[238]^x[236]^x[230]^x[227]^x[213]^x[202]^x[191]^x[190]^x[189]^x[186]^x[184]^x[180]^x[179]^x[178]^x[176]^x[175]^x[174]^x[165]^x[164]^x[163]^x[153]^x[152]^x[142]^x[138]^x[124]^x[122]^x[120]^x[116]^x[115]^x[114]^x[113]^x[110]^x[108]^x[104]^x[102]^x[100]^x[93]^x[88]^x[78]^x[76]^x[72]^x[67]^x[66]^x[59]^x[38]^x[26]^x[16]^x[15]^x[14]^x[5]^x[4]^x[3]^x[0];
	x_new[151]=x[372]^x[366]^x[361]^x[355]^x[345]^x[344]^x[343]^x[342]^x[335]^x[334]^x[331]^x[324]^x[323]^x[322]^x[316]^x[283]^x[281]^x[279]^x[277]^x[274]^x[272]^x[268]^x[266]^x[259]^x[252]^x[247]^x[246]^x[241]^x[240]^x[237]^x[235]^x[229]^x[226]^x[212]^x[201]^x[190]^x[189]^x[188]^x[185]^x[183]^x[179]^x[178]^x[177]^x[175]^x[174]^x[173]^x[164]^x[163]^x[162]^x[152]^x[151]^x[141]^x[137]^x[123]^x[121]^x[119]^x[115]^x[114]^x[113]^x[112]^x[109]^x[107]^x[103]^x[101]^x[99]^x[92]^x[87]^x[77]^x[75]^x[71]^x[66]^x[65]^x[58]^x[25]^x[15]^x[14]^x[13]^x[4]^x[3]^x[2];
	x_new[150]=x[371]^x[365]^x[360]^x[354]^x[344]^x[343]^x[342]^x[341]^x[334]^x[333]^x[330]^x[323]^x[322]^x[321]^x[315]^x[282]^x[280]^x[278]^x[276]^x[273]^x[271]^x[267]^x[265]^x[258]^x[251]^x[246]^x[245]^x[240]^x[239]^x[236]^x[234]^x[228]^x[225]^x[211]^x[200]^x[189]^x[188]^x[187]^x[184]^x[182]^x[178]^x[177]^x[176]^x[174]^x[173]^x[172]^x[163]^x[162]^x[161]^x[151]^x[150]^x[140]^x[136]^x[122]^x[120]^x[118]^x[114]^x[113]^x[112]^x[111]^x[108]^x[106]^x[102]^x[100]^x[98]^x[91]^x[86]^x[76]^x[74]^x[70]^x[65]^x[64]^x[57]^x[24]^x[14]^x[13]^x[12]^x[3]^x[2]^x[1];
	x_new[149]=x[370]^x[364]^x[359]^x[353]^x[343]^x[340]^x[333]^x[332]^x[330]^x[329]^x[322]^x[321]^x[314]^x[281]^x[279]^x[277]^x[275]^x[272]^x[270]^x[267]^x[264]^x[257]^x[256]^x[250]^x[245]^x[244]^x[239]^x[238]^x[235]^x[233]^x[227]^x[224]^x[210]^x[199]^x[188]^x[187]^x[186]^x[183]^x[181]^x[177]^x[176]^x[175]^x[173]^x[172]^x[171]^x[162]^x[161]^x[160]^x[150]^x[149]^x[139]^x[135]^x[121]^x[119]^x[117]^x[113]^x[112]^x[111]^x[110]^x[106]^x[105]^x[100]^x[99]^x[97]^x[96]^x[90]^x[85]^x[75]^x[73]^x[69]^x[64]^x[56]^x[23]^x[13]^x[12]^x[11]^x[2]^x[1]^x[0];
	x_new[148]=x[369]^x[363]^x[358]^x[352]^x[351]^x[350]^x[342]^x[339]^x[332]^x[331]^x[328]^x[321]^x[320]^x[287]^x[286]^x[282]^x[281]^x[278]^x[276]^x[274]^x[270]^x[265]^x[256]^x[255]^x[249]^x[244]^x[243]^x[238]^x[237]^x[232]^x[226]^x[209]^x[198]^x[191]^x[187]^x[186]^x[185]^x[182]^x[180]^x[174]^x[172]^x[171]^x[165]^x[161]^x[160]^x[149]^x[148]^x[138]^x[134]^x[127]^x[126]^x[122]^x[120]^x[118]^x[112]^x[110]^x[106]^x[105]^x[104]^x[100]^x[99]^x[98]^x[96]^x[95]^x[84]^x[83]^x[72]^x[34]^x[31]^x[22]^x[12]^x[11]^x[1]^x[0];
	x_new[147]=x[368]^x[357]^x[351]^x[350]^x[349]^x[341]^x[340]^x[339]^x[338]^x[331]^x[329]^x[327]^x[320]^x[287]^x[285]^x[277]^x[274]^x[273]^x[266]^x[264]^x[263]^x[254]^x[248]^x[243]^x[242]^x[237]^x[236]^x[231]^x[225]^x[208]^x[197]^x[191]^x[190]^x[186]^x[185]^x[184]^x[181]^x[179]^x[175]^x[173]^x[171]^x[160]^x[148]^x[147]^x[137]^x[133]^x[127]^x[125]^x[121]^x[119]^x[117]^x[115]^x[111]^x[109]^x[106]^x[105]^x[104]^x[103]^x[100]^x[99]^x[98]^x[97]^x[94]^x[83]^x[82]^x[71]^x[31]^x[30]^x[21]^x[11]^x[0];
	x_new[146]=x[367]^x[356]^x[351]^x[350]^x[349]^x[348]^x[340]^x[339]^x[338]^x[337]^x[328]^x[326]^x[286]^x[284]^x[276]^x[273]^x[272]^x[265]^x[263]^x[262]^x[253]^x[247]^x[242]^x[241]^x[236]^x[235]^x[230]^x[224]^x[207]^x[196]^x[191]^x[190]^x[189]^x[185]^x[184]^x[183]^x[180]^x[178]^x[174]^x[172]^x[147]^x[146]^x[136]^x[132]^x[126]^x[124]^x[120]^x[118]^x[116]^x[114]^x[110]^x[108]^x[105]^x[104]^x[103]^x[102]^x[99]^x[98]^x[97]^x[96]^x[93]^x[82]^x[81]^x[70]^x[31]^x[30]^x[29]^x[20];
	x_new[145]=x[366]^x[355]^x[350]^x[349]^x[348]^x[347]^x[339]^x[338]^x[337]^x[336]^x[327]^x[325]^x[285]^x[283]^x[278]^x[277]^x[275]^x[266]^x[264]^x[262]^x[260]^x[256]^x[252]^x[246]^x[241]^x[240]^x[235]^x[229]^x[206]^x[195]^x[190]^x[189]^x[188]^x[184]^x[183]^x[182]^x[179]^x[177]^x[173]^x[171]^x[146]^x[145]^x[135]^x[131]^x[125]^x[123]^x[119]^x[118]^x[115]^x[113]^x[109]^x[107]^x[106]^x[104]^x[103]^x[102]^x[101]^x[98]^x[97]^x[92]^x[81]^x[80]^x[69]^x[30]^x[29]^x[28]^x[19];
	x_new[144]=x[365]^x[354]^x[349]^x[348]^x[347]^x[346]^x[338]^x[337]^x[336]^x[335]^x[326]^x[324]^x[284]^x[282]^x[276]^x[274]^x[271]^x[265]^x[263]^x[261]^x[260]^x[259]^x[251]^x[245]^x[240]^x[239]^x[234]^x[228]^x[205]^x[194]^x[189]^x[188]^x[187]^x[183]^x[182]^x[181]^x[178]^x[176]^x[172]^x[170]^x[145]^x[144]^x[134]^x[130]^x[124]^x[122]^x[118]^x[114]^x[112]^x[108]^x[106]^x[105]^x[103]^x[102]^x[101]^x[100]^x[97]^x[96]^x[91]^x[80]^x[79]^x[68]^x[29]^x[28]^x[27]^x[18];
	x_new[143]=x[364]^x[353]^x[348]^x[347]^x[346]^x[345]^x[337]^x[336]^x[335]^x[334]^x[325]^x[323]^x[283]^x[281]^x[277]^x[275]^x[273]^x[271]^x[270]^x[266]^x[264]^x[262]^x[259]^x[258]^x[250]^x[244]^x[239]^x[238]^x[233]^x[227]^x[204]^x[193]^x[188]^x[187]^x[186]^x[182]^x[181]^x[180]^x[177]^x[175]^x[170]^x[169]^x[160]^x[144]^x[143]^x[133]^x[129]^x[123]^x[121]^x[113]^x[111]^x[107]^x[106]^x[105]^x[104]^x[102]^x[101]^x[100]^x[99]^x[96]^x[90]^x[79]^x[78]^x[67]^x[28]^x[27]^x[26]^x[17];
	x_new[142]=x[363]^x[352]^x[347]^x[346]^x[345]^x[344]^x[336]^x[335]^x[334]^x[333]^x[324]^x[322]^x[282]^x[280]^x[276]^x[274]^x[272]^x[270]^x[269]^x[265]^x[263]^x[261]^x[258]^x[257]^x[249]^x[243]^x[238]^x[237]^x[232]^x[226]^x[203]^x[192]^x[187]^x[186]^x[185]^x[181]^x[180]^x[179]^x[176]^x[174]^x[170]^x[169]^x[168]^x[143]^x[142]^x[132]^x[128]^x[122]^x[120]^x[112]^x[110]^x[106]^x[105]^x[104]^x[103]^x[101]^x[100]^x[99]^x[98]^x[89]^x[78]^x[77]^x[66]^x[27]^x[26]^x[25]^x[16];
	x_new[141]=x[346]^x[345]^x[344]^x[343]^x[335]^x[334]^x[333]^x[332]^x[323]^x[321]^x[281]^x[279]^x[275]^x[273]^x[271]^x[269]^x[268]^x[264]^x[262]^x[260]^x[257]^x[256]^x[248]^x[242]^x[237]^x[236]^x[231]^x[225]^x[186]^x[185]^x[184]^x[180]^x[179]^x[178]^x[175]^x[173]^x[169]^x[168]^x[167]^x[142]^x[141]^x[131]^x[121]^x[119]^x[111]^x[109]^x[105]^x[104]^x[103]^x[102]^x[100]^x[99]^x[98]^x[97]^x[88]^x[77]^x[76]^x[65]^x[26]^x[25]^x[24]^x[15];
	x_new[140]=x[345]^x[344]^x[343]^x[342]^x[334]^x[333]^x[332]^x[331]^x[322]^x[320]^x[280]^x[278]^x[274]^x[272]^x[270]^x[268]^x[263]^x[261]^x[259]^x[247]^x[241]^x[236]^x[235]^x[230]^x[224]^x[185]^x[184]^x[183]^x[179]^x[178]^x[177]^x[174]^x[172]^x[168]^x[167]^x[166]^x[141]^x[140]^x[130]^x[120]^x[118]^x[110]^x[108]^x[104]^x[103]^x[102]^x[101]^x[99]^x[98]^x[97]^x[96]^x[87]^x[76]^x[75]^x[64]^x[25]^x[24]^x[23]^x[14];
	x_new[139]=x[344]^x[343]^x[342]^x[333]^x[331]^x[320]^x[279]^x[278]^x[273]^x[272]^x[269]^x[262]^x[261]^x[258]^x[246]^x[240]^x[235]^x[229]^x[184]^x[183]^x[182]^x[178]^x[177]^x[176]^x[173]^x[171]^x[167]^x[166]^x[165]^x[140]^x[139]^x[129]^x[119]^x[118]^x[109]^x[103]^x[102]^x[101]^x[98]^x[97]^x[96]^x[86]^x[75]^x[24]^x[23]^x[22]^x[13];
	x_new[138]=x[343]^x[342]^x[341]^x[332]^x[331]^x[330]^x[320]^x[278]^x[272]^x[268]^x[266]^x[261]^x[257]^x[245]^x[239]^x[234]^x[228]^x[183]^x[182]^x[181]^x[177]^x[176]^x[175]^x[172]^x[170]^x[166]^x[165]^x[164]^x[139]^x[138]^x[128]^x[118]^x[108]^x[106]^x[102]^x[101]^x[100]^x[97]^x[96]^x[85]^x[74]^x[23]^x[22]^x[21]^x[12];
	x_new[137]=x[351]^x[350]^x[342]^x[341]^x[339]^x[331]^x[329]^x[285]^x[277]^x[276]^x[275]^x[267]^x[263]^x[256]^x[244]^x[238]^x[233]^x[227]^x[186]^x[182]^x[181]^x[180]^x[176]^x[175]^x[174]^x[171]^x[169]^x[165]^x[163]^x[159]^x[137]^x[117]^x[116]^x[115]^x[111]^x[110]^x[109]^x[107]^x[105]^x[101]^x[99]^x[96]^x[84]^x[73]^x[22]^x[21]^x[20]^x[11];
	x_new[136]=x[349]^x[341]^x[340]^x[339]^x[338]^x[330]^x[328]^x[287]^x[284]^x[276]^x[275]^x[274]^x[262]^x[243]^x[237]^x[232]^x[226]^x[181]^x[180]^x[179]^x[175]^x[174]^x[173]^x[170]^x[168]^x[164]^x[162]^x[158]^x[136]^x[127]^x[121]^x[116]^x[114]^x[110]^x[108]^x[104]^x[98]^x[83]^x[72]^x[21]^x[20]^x[19]^x[10];
	x_new[135]=x[348]^x[340]^x[339]^x[338]^x[337]^x[329]^x[327]^x[286]^x[283]^x[275]^x[274]^x[273]^x[261]^x[242]^x[236]^x[231]^x[225]^x[180]^x[179]^x[178]^x[174]^x[173]^x[172]^x[169]^x[167]^x[163]^x[161]^x[157]^x[135]^x[126]^x[120]^x[115]^x[113]^x[109]^x[107]^x[103]^x[97]^x[82]^x[71]^x[42]^x[20]^x[19]^x[18]^x[9];
	x_new[134]=x[347]^x[339]^x[338]^x[337]^x[336]^x[328]^x[326]^x[285]^x[282]^x[274]^x[273]^x[272]^x[260]^x[241]^x[235]^x[230]^x[224]^x[179]^x[178]^x[177]^x[173]^x[172]^x[171]^x[168]^x[166]^x[162]^x[160]^x[156]^x[134]^x[125]^x[119]^x[114]^x[112]^x[108]^x[106]^x[102]^x[96]^x[81]^x[70]^x[41]^x[19]^x[18]^x[17]^x[8];
	x_new[133]=x[346]^x[338]^x[337]^x[335]^x[327]^x[309]^x[298]^x[284]^x[281]^x[278]^x[273]^x[271]^x[261]^x[259]^x[256]^x[240]^x[229]^x[182]^x[178]^x[177]^x[176]^x[167]^x[165]^x[160]^x[155]^x[133]^x[124]^x[113]^x[111]^x[107]^x[105]^x[96]^x[80]^x[74]^x[69]^x[68]^x[40]^x[18]^x[17]^x[16]^x[7];
	x_new[132]=x[345]^x[337]^x[336]^x[335]^x[334]^x[326]^x[324]^x[308]^x[297]^x[283]^x[280]^x[277]^x[272]^x[270]^x[266]^x[260]^x[258]^x[239]^x[228]^x[177]^x[176]^x[175]^x[166]^x[164]^x[154]^x[132]^x[123]^x[112]^x[110]^x[104]^x[100]^x[79]^x[73]^x[68]^x[67]^x[39]^x[17]^x[16]^x[15]^x[6];
	x_new[131]=x[344]^x[336]^x[335]^x[334]^x[333]^x[325]^x[323]^x[307]^x[296]^x[282]^x[279]^x[276]^x[271]^x[269]^x[265]^x[259]^x[257]^x[238]^x[227]^x[176]^x[175]^x[174]^x[165]^x[163]^x[153]^x[131]^x[122]^x[111]^x[109]^x[103]^x[99]^x[78]^x[72]^x[67]^x[66]^x[38]^x[16]^x[15]^x[14]^x[5];
	x_new[130]=x[343]^x[335]^x[334]^x[333]^x[332]^x[324]^x[322]^x[306]^x[295]^x[281]^x[278]^x[275]^x[270]^x[268]^x[264]^x[258]^x[256]^x[237]^x[226]^x[175]^x[174]^x[173]^x[164]^x[162]^x[152]^x[130]^x[121]^x[110]^x[108]^x[102]^x[98]^x[77]^x[71]^x[66]^x[65]^x[37]^x[15]^x[14]^x[13]^x[4];
	x_new[129]=x[342]^x[334]^x[333]^x[332]^x[331]^x[323]^x[321]^x[305]^x[294]^x[280]^x[274]^x[269]^x[267]^x[263]^x[257]^x[236]^x[225]^x[174]^x[173]^x[172]^x[163]^x[161]^x[151]^x[129]^x[120]^x[109]^x[107]^x[101]^x[97]^x[76]^x[70]^x[65]^x[64]^x[14]^x[13]^x[12]^x[3];
	x_new[128]=x[342]^x[333]^x[332]^x[331]^x[322]^x[304]^x[293]^x[279]^x[273]^x[268]^x[267]^x[262]^x[235]^x[224]^x[173]^x[172]^x[171]^x[162]^x[160]^x[150]^x[128]^x[119]^x[108]^x[107]^x[101]^x[75]^x[69]^x[64]^x[13]^x[12]^x[11]^x[2];
	x_new[127]=x[375]^x[370]^x[365]^x[362]^x[359]^x[354]^x[352]^x[348]^x[342]^x[337]^x[331]^x[319]^x[318]^x[311]^x[310]^x[309]^x[308]^x[307]^x[299]^x[289]^x[250]^x[249]^x[245]^x[240]^x[238]^x[236]^x[235]^x[234]^x[231]^x[229]^x[225]^x[223]^x[222]^x[217]^x[216]^x[213]^x[211]^x[207]^x[205]^x[202]^x[196]^x[188]^x[177]^x[159]^x[155]^x[154]^x[153]^x[144]^x[135]^x[134]^x[129]^x[127]^x[117]^x[113]^x[107]^x[101]^x[96]^x[90]^x[89]^x[85]^x[84]^x[83]^x[80]^x[79]^x[77]^x[76]^x[75]^x[70]^x[65]^x[64]^x[63]^x[62]^x[53]^x[51]^x[42]^x[2];
	x_new[126]=x[383]^x[374]^x[369]^x[364]^x[362]^x[361]^x[358]^x[353]^x[347]^x[341]^x[336]^x[330]^x[318]^x[317]^x[310]^x[309]^x[308]^x[306]^x[298]^x[297]^x[288]^x[254]^x[253]^x[242]^x[235]^x[234]^x[230]^x[224]^x[222]^x[221]^x[216]^x[215]^x[212]^x[210]^x[206]^x[204]^x[201]^x[195]^x[187]^x[176]^x[158]^x[152]^x[134]^x[133]^x[128]^x[127]^x[126]^x[116]^x[112]^x[100]^x[94]^x[88]^x[82]^x[76]^x[75]^x[74]^x[69]^x[68]^x[64]^x[62]^x[61]^x[52]^x[50]^x[41];
	x_new[125]=x[382]^x[373]^x[368]^x[363]^x[361]^x[360]^x[357]^x[352]^x[346]^x[340]^x[335]^x[329]^x[319]^x[318]^x[317]^x[316]^x[309]^x[308]^x[305]^x[298]^x[297]^x[296]^x[255]^x[253]^x[252]^x[241]^x[233]^x[229]^x[221]^x[220]^x[215]^x[214]^x[211]^x[209]^x[205]^x[203]^x[200]^x[194]^x[186]^x[175]^x[157]^x[151]^x[133]^x[126]^x[125]^x[115]^x[111]^x[99]^x[95]^x[93]^x[89]^x[87]^x[83]^x[81]^x[77]^x[75]^x[73]^x[67]^x[61]^x[60]^x[51]^x[49]^x[40]^x[11]^x[0];
	x_new[124]=x[383]^x[381]^x[372]^x[367]^x[360]^x[359]^x[356]^x[345]^x[339]^x[334]^x[328]^x[318]^x[317]^x[316]^x[315]^x[308]^x[307]^x[304]^x[297]^x[296]^x[295]^x[254]^x[252]^x[251]^x[240]^x[232]^x[228]^x[220]^x[219]^x[214]^x[213]^x[210]^x[208]^x[204]^x[202]^x[199]^x[193]^x[185]^x[174]^x[156]^x[150]^x[132]^x[125]^x[124]^x[114]^x[110]^x[98]^x[94]^x[92]^x[88]^x[86]^x[82]^x[80]^x[76]^x[74]^x[72]^x[66]^x[60]^x[59]^x[50]^x[48]^x[39]^x[10];
	x_new[123]=x[382]^x[380]^x[371]^x[366]^x[359]^x[358]^x[355]^x[344]^x[338]^x[333]^x[327]^x[317]^x[316]^x[315]^x[314]^x[307]^x[306]^x[303]^x[296]^x[295]^x[294]^x[253]^x[251]^x[250]^x[239]^x[231]^x[227]^x[219]^x[218]^x[213]^x[212]^x[209]^x[207]^x[203]^x[201]^x[198]^x[192]^x[184]^x[173]^x[155]^x[149]^x[131]^x[124]^x[123]^x[113]^x[109]^x[97]^x[93]^x[91]^x[87]^x[85]^x[81]^x[79]^x[75]^x[73]^x[71]^x[65]^x[59]^x[58]^x[49]^x[47]^x[38]^x[9];
	x_new[122]=x[381]^x[379]^x[370]^x[365]^x[358]^x[357]^x[354]^x[343]^x[337]^x[332]^x[326]^x[316]^x[315]^x[313]^x[306]^x[305]^x[302]^x[295]^x[294]^x[293]^x[287]^x[255]^x[254]^x[252]^x[248]^x[245]^x[244]^x[243]^x[239]^x[237]^x[235]^x[230]^x[226]^x[224]^x[223]^x[218]^x[217]^x[212]^x[211]^x[208]^x[206]^x[200]^x[197]^x[183]^x[172]^x[159]^x[154]^x[150]^x[149]^x[148]^x[139]^x[138]^x[130]^x[123]^x[122]^x[112]^x[108]^x[96]^x[95]^x[94]^x[92]^x[86]^x[85]^x[84]^x[83]^x[80]^x[78]^x[75]^x[74]^x[72]^x[70]^x[69]^x[63]^x[58]^x[48]^x[46]^x[42]^x[37]^x[36]^x[29];
	x_new[121]=x[380]^x[378]^x[369]^x[364]^x[357]^x[356]^x[353]^x[342]^x[336]^x[331]^x[325]^x[315]^x[314]^x[313]^x[312]^x[305]^x[304]^x[301]^x[294]^x[293]^x[292]^x[286]^x[253]^x[251]^x[249]^x[248]^x[247]^x[244]^x[242]^x[238]^x[237]^x[236]^x[229]^x[225]^x[222]^x[217]^x[216]^x[211]^x[210]^x[207]^x[205]^x[199]^x[196]^x[182]^x[171]^x[159]^x[158]^x[153]^x[148]^x[147]^x[138]^x[137]^x[129]^x[122]^x[121]^x[111]^x[107]^x[93]^x[91]^x[89]^x[85]^x[84]^x[83]^x[82]^x[79]^x[77]^x[73]^x[71]^x[69]^x[62]^x[57]^x[47]^x[45]^x[41]^x[36]^x[35]^x[28]^x[7];
	x_new[120]=x[379]^x[377]^x[368]^x[363]^x[356]^x[355]^x[352]^x[341]^x[335]^x[330]^x[324]^x[314]^x[313]^x[312]^x[311]^x[304]^x[303]^x[300]^x[293]^x[292]^x[291]^x[285]^x[252]^x[250]^x[248]^x[247]^x[246]^x[243]^x[241]^x[237]^x[236]^x[235]^x[228]^x[224]^x[221]^x[216]^x[215]^x[210]^x[209]^x[206]^x[204]^x[198]^x[195]^x[181]^x[170]^x[159]^x[158]^x[157]^x[152]^x[147]^x[146]^x[138]^x[137]^x[136]^x[128]^x[121]^x[120]^x[110]^x[106]^x[92]^x[90]^x[88]^x[84]^x[83]^x[82]^x[81]^x[78]^x[76]^x[72]^x[70]^x[68]^x[61]^x[56]^x[46]^x[44]^x[40]^x[35]^x[34]^x[27]^x[6];
	x_new[119]=x[378]^x[376]^x[367]^x[355]^x[354]^x[340]^x[334]^x[329]^x[323]^x[313]^x[312]^x[311]^x[310]^x[303]^x[302]^x[299]^x[292]^x[291]^x[290]^x[284]^x[251]^x[249]^x[247]^x[245]^x[242]^x[240]^x[236]^x[234]^x[227]^x[220]^x[215]^x[214]^x[209]^x[208]^x[205]^x[203]^x[197]^x[194]^x[180]^x[169]^x[158]^x[157]^x[156]^x[151]^x[146]^x[145]^x[137]^x[136]^x[135]^x[120]^x[119]^x[109]^x[105]^x[91]^x[89]^x[87]^x[83]^x[82]^x[81]^x[80]^x[77]^x[75]^x[71]^x[69]^x[67]^x[60]^x[55]^x[45]^x[43]^x[39]^x[34]^x[33]^x[26];
	x_new[118]=x[377]^x[375]^x[366]^x[354]^x[353]^x[339]^x[333]^x[328]^x[322]^x[312]^x[311]^x[310]^x[309]^x[302]^x[301]^x[298]^x[291]^x[290]^x[289]^x[283]^x[250]^x[248]^x[246]^x[244]^x[241]^x[239]^x[235]^x[233]^x[226]^x[219]^x[214]^x[213]^x[208]^x[207]^x[204]^x[202]^x[196]^x[193]^x[179]^x[168]^x[157]^x[156]^x[155]^x[150]^x[145]^x[144]^x[136]^x[135]^x[134]^x[119]^x[118]^x[108]^x[104]^x[90]^x[88]^x[86]^x[82]^x[81]^x[80]^x[79]^x[76]^x[74]^x[70]^x[68]^x[66]^x[59]^x[54]^x[44]^x[42]^x[38]^x[33]^x[32]^x[25];
	x_new[117]=x[376]^x[374]^x[365]^x[353]^x[352]^x[338]^x[332]^x[327]^x[321]^x[311]^x[308]^x[301]^x[300]^x[298]^x[297]^x[290]^x[289]^x[282]^x[249]^x[247]^x[245]^x[243]^x[240]^x[238]^x[235]^x[232]^x[225]^x[224]^x[218]^x[213]^x[212]^x[207]^x[206]^x[203]^x[201]^x[195]^x[192]^x[178]^x[167]^x[156]^x[155]^x[154]^x[149]^x[144]^x[143]^x[135]^x[134]^x[133]^x[118]^x[117]^x[107]^x[103]^x[89]^x[87]^x[85]^x[81]^x[80]^x[79]^x[78]^x[74]^x[73]^x[68]^x[67]^x[65]^x[64]^x[58]^x[53]^x[43]^x[41]^x[37]^x[32]^x[24];
	x_new[116]=x[383]^x[375]^x[373]^x[364]^x[362]^x[352]^x[337]^x[331]^x[326]^x[320]^x[319]^x[318]^x[310]^x[307]^x[300]^x[299]^x[296]^x[289]^x[288]^x[255]^x[254]^x[250]^x[249]^x[246]^x[244]^x[242]^x[238]^x[233]^x[224]^x[223]^x[217]^x[212]^x[211]^x[206]^x[205]^x[200]^x[194]^x[177]^x[166]^x[155]^x[154]^x[148]^x[144]^x[142]^x[134]^x[117]^x[116]^x[106]^x[102]^x[95]^x[94]^x[90]^x[88]^x[86]^x[80]^x[78]^x[74]^x[73]^x[72]^x[68]^x[67]^x[66]^x[64]^x[63]^x[52]^x[51]^x[40]^x[2];
	x_new[115]=x[383]^x[382]^x[374]^x[372]^x[363]^x[362]^x[361]^x[336]^x[325]^x[319]^x[318]^x[317]^x[309]^x[308]^x[307]^x[306]^x[299]^x[297]^x[295]^x[288]^x[255]^x[253]^x[245]^x[242]^x[241]^x[234]^x[232]^x[231]^x[222]^x[216]^x[211]^x[210]^x[205]^x[204]^x[199]^x[193]^x[176]^x[165]^x[154]^x[147]^x[141]^x[133]^x[116]^x[115]^x[105]^x[101]^x[95]^x[93]^x[89]^x[87]^x[85]^x[83]^x[79]^x[77]^x[74]^x[73]^x[72]^x[71]^x[68]^x[67]^x[66]^x[65]^x[62]^x[51]^x[50]^x[39];
	x_new[114]=x[382]^x[381]^x[373]^x[371]^x[362]^x[361]^x[360]^x[335]^x[324]^x[319]^x[318]^x[317]^x[316]^x[308]^x[307]^x[306]^x[305]^x[296]^x[294]^x[254]^x[252]^x[244]^x[241]^x[240]^x[233]^x[231]^x[230]^x[221]^x[215]^x[210]^x[209]^x[204]^x[203]^x[198]^x[192]^x[175]^x[164]^x[146]^x[140]^x[115]^x[114]^x[104]^x[100]^x[94]^x[92]^x[88]^x[86]^x[84]^x[82]^x[78]^x[76]^x[73]^x[72]^x[71]^x[70]^x[67]^x[66]^x[65]^x[64]^x[61]^x[50]^x[49]^x[38];
	x_new[113]=x[381]^x[380]^x[372]^x[370]^x[361]^x[360]^x[359]^x[334]^x[323]^x[318]^x[317]^x[316]^x[315]^x[307]^x[306]^x[305]^x[304]^x[295]^x[293]^x[253]^x[251]^x[246]^x[245]^x[243]^x[234]^x[232]^x[230]^x[228]^x[224]^x[220]^x[214]^x[209]^x[208]^x[203]^x[197]^x[174]^x[163]^x[145]^x[139]^x[114]^x[113]^x[103]^x[99]^x[93]^x[91]^x[87]^x[86]^x[83]^x[81]^x[77]^x[75]^x[74]^x[72]^x[71]^x[70]^x[69]^x[66]^x[65]^x[60]^x[49]^x[48]^x[37];
	x_new[112]=x[380]^x[379]^x[371]^x[369]^x[360]^x[359]^x[358]^x[333]^x[322]^x[317]^x[316]^x[315]^x[314]^x[306]^x[305]^x[304]^x[303]^x[294]^x[292]^x[252]^x[250]^x[244]^x[242]^x[239]^x[233]^x[231]^x[229]^x[228]^x[227]^x[219]^x[213]^x[208]^x[207]^x[202]^x[196]^x[173]^x[162]^x[144]^x[138]^x[113]^x[112]^x[102]^x[98]^x[92]^x[90]^x[86]^x[82]^x[80]^x[76]^x[74]^x[73]^x[71]^x[70]^x[69]^x[68]^x[65]^x[64]^x[59]^x[48]^x[47]^x[36];
	x_new[111]=x[379]^x[378]^x[370]^x[368]^x[359]^x[358]^x[357]^x[332]^x[321]^x[316]^x[315]^x[314]^x[313]^x[305]^x[304]^x[303]^x[302]^x[293]^x[291]^x[251]^x[249]^x[245]^x[243]^x[241]^x[239]^x[238]^x[234]^x[232]^x[230]^x[227]^x[226]^x[218]^x[212]^x[207]^x[206]^x[201]^x[195]^x[172]^x[161]^x[143]^x[139]^x[138]^x[137]^x[128]^x[112]^x[111]^x[101]^x[97]^x[91]^x[89]^x[81]^x[79]^x[75]^x[74]^x[73]^x[72]^x[70]^x[69]^x[68]^x[67]^x[64]^x[58]^x[47]^x[46]^x[35];
	x_new[110]=x[378]^x[377]^x[369]^x[367]^x[358]^x[357]^x[356]^x[331]^x[320]^x[315]^x[314]^x[313]^x[312]^x[304]^x[303]^x[302]^x[301]^x[292]^x[290]^x[250]^x[248]^x[244]^x[242]^x[240]^x[238]^x[237]^x[233]^x[231]^x[229]^x[226]^x[225]^x[217]^x[211]^x[206]^x[205]^x[200]^x[194]^x[171]^x[160]^x[142]^x[137]^x[136]^x[111]^x[110]^x[100]^x[96]^x[90]^x[88]^x[80]^x[78]^x[74]^x[73]^x[72]^x[71]^x[69]^x[68]^x[67]^x[66]^x[57]^x[46]^x[45]^x[34];
	x_new[109]=x[377]^x[376]^x[368]^x[366]^x[357]^x[356]^x[355]^x[314]^x[313]^x[312]^x[311]^x[303]^x[302]^x[301]^x[300]^x[291]^x[289]^x[249]^x[247]^x[243]^x[241]^x[239]^x[237]^x[236]^x[232]^x[230]^x[228]^x[225]^x[224]^x[216]^x[210]^x[205]^x[204]^x[199]^x[193]^x[141]^x[136]^x[135]^x[110]^x[109]^x[99]^x[89]^x[87]^x[79]^x[77]^x[73]^x[72]^x[71]^x[70]^x[68]^x[67]^x[66]^x[65]^x[56]^x[45]^x[44]^x[33];
	x_new[108]=x[376]^x[375]^x[367]^x[365]^x[356]^x[355]^x[354]^x[313]^x[312]^x[311]^x[310]^x[302]^x[301]^x[300]^x[299]^x[290]^x[288]^x[248]^x[246]^x[242]^x[240]^x[238]^x[236]^x[231]^x[229]^x[227]^x[215]^x[209]^x[204]^x[203]^x[198]^x[192]^x[140]^x[135]^x[134]^x[109]^x[108]^x[98]^x[88]^x[86]^x[78]^x[76]^x[72]^x[71]^x[70]^x[69]^x[67]^x[66]^x[65]^x[64]^x[55]^x[44]^x[43]^x[32];
	x_new[107]=x[375]^x[374]^x[366]^x[364]^x[355]^x[354]^x[353]^x[312]^x[311]^x[310]^x[301]^x[299]^x[288]^x[247]^x[246]^x[241]^x[240]^x[237]^x[230]^x[229]^x[226]^x[214]^x[208]^x[203]^x[197]^x[139]^x[134]^x[133]^x[108]^x[107]^x[97]^x[87]^x[86]^x[77]^x[71]^x[70]^x[69]^x[66]^x[65]^x[64]^x[54]^x[43];
	x_new[106]=x[374]^x[373]^x[365]^x[363]^x[354]^x[353]^x[352]^x[311]^x[310]^x[309]^x[300]^x[299]^x[298]^x[288]^x[246]^x[240]^x[236]^x[234]^x[229]^x[225]^x[213]^x[207]^x[202]^x[196]^x[138]^x[133]^x[132]^x[107]^x[106]^x[96]^x[86]^x[76]^x[74]^x[70]^x[69]^x[68]^x[65]^x[64]^x[53]^x[42];
	x_new[105]=x[383]^x[373]^x[372]^x[364]^x[353]^x[352]^x[319]^x[318]^x[310]^x[309]^x[307]^x[299]^x[297]^x[253]^x[245]^x[244]^x[243]^x[235]^x[231]^x[224]^x[212]^x[206]^x[201]^x[195]^x[154]^x[137]^x[131]^x[127]^x[105]^x[85]^x[84]^x[83]^x[79]^x[78]^x[77]^x[75]^x[73]^x[69]^x[67]^x[64]^x[52]^x[41];
	x_new[104]=x[383]^x[382]^x[372]^x[371]^x[363]^x[362]^x[352]^x[317]^x[309]^x[308]^x[307]^x[306]^x[298]^x[296]^x[255]^x[252]^x[244]^x[243]^x[242]^x[230]^x[211]^x[205]^x[200]^x[194]^x[136]^x[130]^x[126]^x[104]^x[95]^x[89]^x[84]^x[82]^x[78]^x[76]^x[72]^x[66]^x[51]^x[40];
	x_new[103]=x[383]^x[382]^x[381]^x[371]^x[370]^x[361]^x[316]^x[308]^x[307]^x[306]^x[305]^x[297]^x[295]^x[254]^x[251]^x[243]^x[242]^x[241]^x[229]^x[210]^x[204]^x[199]^x[193]^x[135]^x[129]^x[125]^x[103]^x[94]^x[88]^x[83]^x[81]^x[77]^x[75]^x[71]^x[65]^x[50]^x[39]^x[10];
	x_new[102]=x[382]^x[381]^x[380]^x[370]^x[369]^x[360]^x[315]^x[307]^x[306]^x[305]^x[304]^x[296]^x[294]^x[253]^x[250]^x[242]^x[241]^x[240]^x[228]^x[209]^x[203]^x[198]^x[192]^x[134]^x[128]^x[124]^x[102]^x[93]^x[87]^x[82]^x[80]^x[76]^x[74]^x[70]^x[64]^x[49]^x[38]^x[9];
	x_new[101]=x[381]^x[380]^x[379]^x[369]^x[368]^x[359]^x[314]^x[306]^x[305]^x[303]^x[295]^x[277]^x[266]^x[252]^x[249]^x[246]^x[241]^x[239]^x[229]^x[227]^x[224]^x[208]^x[197]^x[150]^x[140]^x[139]^x[138]^x[133]^x[129]^x[128]^x[123]^x[101]^x[92]^x[81]^x[79]^x[75]^x[73]^x[64]^x[48]^x[42]^x[37]^x[36]^x[8];
	x_new[100]=x[380]^x[379]^x[378]^x[368]^x[367]^x[358]^x[313]^x[305]^x[304]^x[303]^x[302]^x[294]^x[292]^x[276]^x[265]^x[251]^x[248]^x[245]^x[240]^x[238]^x[234]^x[228]^x[226]^x[207]^x[196]^x[139]^x[138]^x[137]^x[132]^x[128]^x[122]^x[100]^x[91]^x[80]^x[78]^x[72]^x[68]^x[47]^x[41]^x[36]^x[35]^x[7];
	x_new[99]=x[379]^x[378]^x[377]^x[367]^x[366]^x[357]^x[312]^x[304]^x[303]^x[302]^x[301]^x[293]^x[291]^x[275]^x[264]^x[250]^x[247]^x[244]^x[239]^x[237]^x[233]^x[227]^x[225]^x[206]^x[195]^x[138]^x[137]^x[136]^x[131]^x[121]^x[99]^x[90]^x[79]^x[77]^x[71]^x[67]^x[46]^x[40]^x[35]^x[34]^x[6];
	x_new[98]=x[378]^x[377]^x[376]^x[366]^x[365]^x[356]^x[311]^x[303]^x[302]^x[301]^x[300]^x[292]^x[290]^x[274]^x[263]^x[249]^x[246]^x[243]^x[238]^x[236]^x[232]^x[226]^x[224]^x[205]^x[194]^x[137]^x[136]^x[135]^x[130]^x[120]^x[98]^x[89]^x[78]^x[76]^x[70]^x[66]^x[45]^x[39]^x[34]^x[33]^x[5];
	x_new[97]=x[377]^x[376]^x[375]^x[365]^x[364]^x[355]^x[310]^x[302]^x[301]^x[300]^x[299]^x[291]^x[289]^x[273]^x[262]^x[248]^x[242]^x[237]^x[235]^x[231]^x[225]^x[204]^x[193]^x[136]^x[135]^x[134]^x[129]^x[119]^x[97]^x[88]^x[77]^x[75]^x[69]^x[65]^x[44]^x[38]^x[33]^x[32];
	x_new[96]=x[376]^x[375]^x[374]^x[364]^x[363]^x[354]^x[310]^x[301]^x[300]^x[299]^x[290]^x[272]^x[261]^x[247]^x[241]^x[236]^x[235]^x[230]^x[203]^x[192]^x[135]^x[134]^x[133]^x[128]^x[118]^x[96]^x[87]^x[76]^x[75]^x[69]^x[43]^x[37]^x[32];
	x_new[95]=x[365]^x[354]^x[343]^x[338]^x[333]^x[330]^x[327]^x[322]^x[320]^x[316]^x[310]^x[305]^x[299]^x[287]^x[286]^x[279]^x[278]^x[277]^x[276]^x[275]^x[267]^x[257]^x[218]^x[217]^x[213]^x[208]^x[206]^x[204]^x[203]^x[202]^x[199]^x[197]^x[193]^x[191]^x[190]^x[185]^x[184]^x[181]^x[179]^x[175]^x[173]^x[170]^x[164]^x[156]^x[145]^x[130]^x[127]^x[123]^x[122]^x[121]^x[112]^x[103]^x[102]^x[97]^x[95]^x[85]^x[81]^x[75]^x[69]^x[64]^x[58]^x[57]^x[53]^x[52]^x[51]^x[48]^x[47]^x[45]^x[44]^x[43]^x[38]^x[33]^x[32]^x[31]^x[30]^x[21]^x[19]^x[10];
	x_new[94]=x[351]^x[342]^x[337]^x[332]^x[330]^x[329]^x[326]^x[321]^x[315]^x[309]^x[304]^x[298]^x[286]^x[285]^x[278]^x[277]^x[276]^x[274]^x[266]^x[265]^x[256]^x[222]^x[221]^x[210]^x[203]^x[202]^x[198]^x[192]^x[190]^x[189]^x[184]^x[183]^x[180]^x[178]^x[174]^x[172]^x[169]^x[163]^x[155]^x[144]^x[126]^x[120]^x[102]^x[101]^x[96]^x[95]^x[94]^x[84]^x[80]^x[68]^x[62]^x[56]^x[50]^x[44]^x[43]^x[42]^x[37]^x[36]^x[32]^x[30]^x[29]^x[20]^x[18]^x[9];
	x_new[93]=x[374]^x[352]^x[350]^x[341]^x[336]^x[331]^x[329]^x[328]^x[325]^x[320]^x[314]^x[308]^x[303]^x[297]^x[287]^x[286]^x[285]^x[284]^x[277]^x[276]^x[273]^x[266]^x[265]^x[264]^x[223]^x[221]^x[220]^x[209]^x[201]^x[197]^x[189]^x[188]^x[183]^x[182]^x[179]^x[177]^x[173]^x[171]^x[168]^x[162]^x[154]^x[143]^x[139]^x[133]^x[128]^x[125]^x[119]^x[101]^x[94]^x[93]^x[83]^x[79]^x[67]^x[63]^x[61]^x[57]^x[55]^x[51]^x[49]^x[45]^x[43]^x[41]^x[35]^x[29]^x[28]^x[19]^x[17]^x[8];
	x_new[92]=x[373]^x[362]^x[351]^x[349]^x[340]^x[335]^x[328]^x[327]^x[324]^x[313]^x[307]^x[302]^x[296]^x[286]^x[285]^x[284]^x[283]^x[276]^x[275]^x[272]^x[265]^x[264]^x[263]^x[222]^x[220]^x[219]^x[208]^x[200]^x[196]^x[188]^x[187]^x[182]^x[181]^x[178]^x[176]^x[172]^x[170]^x[167]^x[161]^x[153]^x[142]^x[138]^x[132]^x[124]^x[118]^x[100]^x[93]^x[92]^x[82]^x[78]^x[66]^x[62]^x[60]^x[56]^x[54]^x[50]^x[48]^x[44]^x[42]^x[40]^x[34]^x[28]^x[27]^x[18]^x[16]^x[7];
	x_new[91]=x[372]^x[361]^x[350]^x[348]^x[339]^x[334]^x[327]^x[326]^x[323]^x[312]^x[306]^x[301]^x[295]^x[285]^x[284]^x[283]^x[282]^x[275]^x[274]^x[271]^x[264]^x[263]^x[262]^x[221]^x[219]^x[218]^x[207]^x[199]^x[195]^x[187]^x[186]^x[181]^x[180]^x[177]^x[175]^x[171]^x[169]^x[166]^x[160]^x[152]^x[141]^x[137]^x[131]^x[123]^x[117]^x[99]^x[92]^x[91]^x[81]^x[77]^x[65]^x[61]^x[59]^x[55]^x[53]^x[49]^x[47]^x[43]^x[41]^x[39]^x[33]^x[27]^x[26]^x[17]^x[15]^x[6];
	x_new[90]=x[381]^x[371]^x[360]^x[349]^x[347]^x[338]^x[333]^x[326]^x[325]^x[322]^x[311]^x[305]^x[300]^x[294]^x[284]^x[283]^x[281]^x[274]^x[273]^x[270]^x[263]^x[262]^x[261]^x[255]^x[223]^x[222]^x[220]^x[216]^x[213]^x[212]^x[211]^x[207]^x[205]^x[203]^x[198]^x[194]^x[192]^x[191]^x[186]^x[185]^x[180]^x[179]^x[176]^x[174]^x[168]^x[165]^x[157]^x[140]^x[127]^x[122]^x[118]^x[117]^x[116]^x[107]^x[106]^x[98]^x[91]^x[90]^x[80]^x[76]^x[64]^x[63]^x[62]^x[60]^x[54]^x[53]^x[52]^x[51]^x[48]^x[46]^x[43]^x[42]^x[40]^x[38]^x[37]^x[31]^x[26]^x[16]^x[14]^x[10]^x[5]^x[4];
	x_new[89]=x[380]^x[348]^x[346]^x[337]^x[332]^x[325]^x[324]^x[321]^x[310]^x[304]^x[299]^x[293]^x[283]^x[282]^x[281]^x[280]^x[273]^x[272]^x[269]^x[262]^x[261]^x[260]^x[254]^x[221]^x[219]^x[217]^x[216]^x[215]^x[212]^x[210]^x[206]^x[205]^x[204]^x[197]^x[193]^x[190]^x[185]^x[184]^x[179]^x[178]^x[175]^x[173]^x[167]^x[164]^x[156]^x[139]^x[135]^x[129]^x[127]^x[126]^x[121]^x[116]^x[115]^x[106]^x[105]^x[97]^x[90]^x[89]^x[79]^x[75]^x[61]^x[59]^x[57]^x[53]^x[52]^x[51]^x[50]^x[47]^x[45]^x[41]^x[39]^x[37]^x[30]^x[25]^x[15]^x[13]^x[9]^x[4]^x[3];
	x_new[88]=x[379]^x[347]^x[345]^x[336]^x[331]^x[324]^x[323]^x[320]^x[309]^x[303]^x[298]^x[292]^x[282]^x[281]^x[280]^x[279]^x[272]^x[271]^x[268]^x[261]^x[260]^x[259]^x[253]^x[220]^x[218]^x[216]^x[215]^x[214]^x[211]^x[209]^x[205]^x[204]^x[203]^x[196]^x[192]^x[189]^x[184]^x[183]^x[178]^x[177]^x[174]^x[172]^x[166]^x[163]^x[155]^x[138]^x[134]^x[128]^x[127]^x[126]^x[125]^x[120]^x[115]^x[114]^x[106]^x[105]^x[104]^x[96]^x[89]^x[88]^x[78]^x[74]^x[60]^x[58]^x[56]^x[52]^x[51]^x[50]^x[49]^x[46]^x[44]^x[40]^x[38]^x[36]^x[29]^x[24]^x[14]^x[12]^x[8]^x[3]^x[2];
	x_new[87]=x[378]^x[368]^x[357]^x[346]^x[344]^x[335]^x[323]^x[322]^x[308]^x[302]^x[297]^x[291]^x[281]^x[280]^x[279]^x[278]^x[271]^x[270]^x[267]^x[260]^x[259]^x[258]^x[252]^x[219]^x[217]^x[215]^x[213]^x[210]^x[208]^x[204]^x[202]^x[195]^x[188]^x[183]^x[182]^x[177]^x[176]^x[173]^x[171]^x[165]^x[162]^x[154]^x[137]^x[126]^x[125]^x[124]^x[119]^x[114]^x[113]^x[105]^x[104]^x[103]^x[88]^x[87]^x[77]^x[73]^x[59]^x[57]^x[55]^x[51]^x[50]^x[49]^x[48]^x[45]^x[43]^x[39]^x[37]^x[35]^x[28]^x[23]^x[13]^x[11]^x[7]^x[2]^x[1];
	x_new[86]=x[377]^x[367]^x[356]^x[345]^x[343]^x[334]^x[322]^x[321]^x[307]^x[301]^x[296]^x[290]^x[280]^x[279]^x[278]^x[277]^x[270]^x[269]^x[266]^x[259]^x[258]^x[257]^x[251]^x[218]^x[216]^x[214]^x[212]^x[209]^x[207]^x[203]^x[201]^x[194]^x[187]^x[182]^x[181]^x[176]^x[175]^x[172]^x[170]^x[164]^x[161]^x[153]^x[136]^x[125]^x[124]^x[123]^x[118]^x[113]^x[112]^x[104]^x[103]^x[102]^x[87]^x[86]^x[76]^x[72]^x[58]^x[56]^x[54]^x[50]^x[49]^x[48]^x[47]^x[44]^x[42]^x[38]^x[36]^x[34]^x[27]^x[22]^x[12]^x[10]^x[6]^x[1]^x[0];
	x_new[85]=x[376]^x[366]^x[355]^x[344]^x[342]^x[333]^x[321]^x[320]^x[306]^x[300]^x[295]^x[289]^x[279]^x[276]^x[269]^x[268]^x[266]^x[265]^x[258]^x[257]^x[250]^x[217]^x[215]^x[213]^x[211]^x[208]^x[206]^x[203]^x[200]^x[193]^x[192]^x[186]^x[181]^x[180]^x[175]^x[174]^x[171]^x[169]^x[163]^x[160]^x[152]^x[135]^x[124]^x[123]^x[122]^x[117]^x[112]^x[111]^x[103]^x[102]^x[101]^x[86]^x[85]^x[75]^x[71]^x[57]^x[55]^x[53]^x[49]^x[48]^x[47]^x[46]^x[42]^x[41]^x[36]^x[35]^x[33]^x[32]^x[26]^x[21]^x[11]^x[9]^x[5]^x[0];
	x_new[84]=x[365]^x[354]^x[351]^x[343]^x[341]^x[332]^x[330]^x[320]^x[305]^x[299]^x[294]^x[288]^x[287]^x[286]^x[278]^x[275]^x[268]^x[267]^x[264]^x[257]^x[256]^x[223]^x[222]^x[218]^x[217]^x[214]^x[212]^x[210]^x[206]^x[201]^x[192]^x[191]^x[185]^x[180]^x[179]^x[174]^x[173]^x[168]^x[162]^x[145]^x[134]^x[130]^x[123]^x[122]^x[116]^x[112]^x[110]^x[102]^x[85]^x[84]^x[74]^x[70]^x[63]^x[62]^x[58]^x[56]^x[54]^x[48]^x[46]^x[42]^x[41]^x[40]^x[36]^x[35]^x[34]^x[32]^x[31]^x[20]^x[19]^x[8];
	x_new[83]=x[351]^x[350]^x[342]^x[340]^x[331]^x[330]^x[329]^x[304]^x[293]^x[287]^x[286]^x[285]^x[277]^x[276]^x[275]^x[274]^x[267]^x[265]^x[263]^x[256]^x[223]^x[221]^x[213]^x[210]^x[209]^x[202]^x[200]^x[199]^x[190]^x[184]^x[179]^x[178]^x[173]^x[172]^x[167]^x[161]^x[144]^x[133]^x[122]^x[115]^x[109]^x[101]^x[84]^x[83]^x[73]^x[69]^x[63]^x[61]^x[57]^x[55]^x[53]^x[51]^x[47]^x[45]^x[42]^x[41]^x[40]^x[39]^x[36]^x[35]^x[34]^x[33]^x[30]^x[19]^x[18]^x[7];
	x_new[82]=x[350]^x[349]^x[341]^x[339]^x[330]^x[329]^x[328]^x[303]^x[292]^x[287]^x[286]^x[285]^x[284]^x[276]^x[275]^x[274]^x[273]^x[264]^x[262]^x[222]^x[220]^x[212]^x[209]^x[208]^x[201]^x[199]^x[198]^x[189]^x[183]^x[178]^x[177]^x[172]^x[171]^x[166]^x[160]^x[143]^x[132]^x[114]^x[108]^x[83]^x[82]^x[72]^x[68]^x[62]^x[60]^x[56]^x[54]^x[52]^x[50]^x[46]^x[44]^x[41]^x[40]^x[39]^x[38]^x[35]^x[34]^x[33]^x[32]^x[29]^x[18]^x[17]^x[6];
	x_new[81]=x[349]^x[348]^x[340]^x[338]^x[329]^x[328]^x[327]^x[302]^x[291]^x[286]^x[285]^x[284]^x[283]^x[275]^x[274]^x[273]^x[272]^x[263]^x[261]^x[221]^x[219]^x[214]^x[213]^x[211]^x[202]^x[200]^x[198]^x[196]^x[192]^x[188]^x[182]^x[177]^x[176]^x[171]^x[165]^x[142]^x[131]^x[113]^x[107]^x[82]^x[81]^x[71]^x[67]^x[61]^x[59]^x[55]^x[54]^x[51]^x[49]^x[45]^x[43]^x[42]^x[40]^x[39]^x[38]^x[37]^x[34]^x[33]^x[28]^x[17]^x[16]^x[5];
	x_new[80]=x[348]^x[347]^x[339]^x[337]^x[328]^x[327]^x[326]^x[301]^x[290]^x[285]^x[284]^x[283]^x[282]^x[274]^x[273]^x[272]^x[271]^x[262]^x[260]^x[220]^x[218]^x[212]^x[210]^x[207]^x[201]^x[199]^x[197]^x[196]^x[195]^x[187]^x[181]^x[176]^x[175]^x[170]^x[164]^x[141]^x[130]^x[112]^x[106]^x[81]^x[80]^x[70]^x[66]^x[60]^x[58]^x[54]^x[50]^x[48]^x[44]^x[42]^x[41]^x[39]^x[38]^x[37]^x[36]^x[33]^x[32]^x[27]^x[16]^x[15]^x[4];
	x_new[79]=x[347]^x[346]^x[338]^x[336]^x[327]^x[326]^x[325]^x[300]^x[289]^x[284]^x[283]^x[282]^x[281]^x[273]^x[272]^x[271]^x[270]^x[261]^x[259]^x[219]^x[217]^x[213]^x[211]^x[209]^x[207]^x[206]^x[202]^x[200]^x[198]^x[195]^x[194]^x[186]^x[180]^x[175]^x[174]^x[169]^x[163]^x[140]^x[129]^x[111]^x[107]^x[106]^x[105]^x[96]^x[80]^x[79]^x[69]^x[65]^x[59]^x[57]^x[49]^x[47]^x[43]^x[42]^x[41]^x[40]^x[38]^x[37]^x[36]^x[35]^x[32]^x[26]^x[15]^x[14]^x[3];
	x_new[78]=x[346]^x[345]^x[337]^x[335]^x[326]^x[325]^x[324]^x[299]^x[288]^x[283]^x[282]^x[281]^x[280]^x[272]^x[271]^x[270]^x[269]^x[260]^x[258]^x[218]^x[216]^x[212]^x[210]^x[208]^x[206]^x[205]^x[201]^x[199]^x[197]^x[194]^x[193]^x[185]^x[179]^x[174]^x[173]^x[168]^x[162]^x[139]^x[128]^x[110]^x[105]^x[104]^x[79]^x[78]^x[68]^x[64]^x[58]^x[56]^x[48]^x[46]^x[42]^x[41]^x[40]^x[39]^x[37]^x[36]^x[35]^x[34]^x[25]^x[14]^x[13]^x[2];
	x_new[77]=x[345]^x[344]^x[336]^x[334]^x[325]^x[324]^x[323]^x[282]^x[281]^x[280]^x[279]^x[271]^x[270]^x[269]^x[268]^x[259]^x[257]^x[217]^x[215]^x[211]^x[209]^x[207]^x[205]^x[204]^x[200]^x[198]^x[196]^x[193]^x[192]^x[184]^x[178]^x[173]^x[172]^x[167]^x[161]^x[109]^x[104]^x[103]^x[78]^x[77]^x[67]^x[57]^x[55]^x[47]^x[45]^x[41]^x[40]^x[39]^x[38]^x[36]^x[35]^x[34]^x[33]^x[24]^x[13]^x[12]^x[1];
	x_new[76]=x[344]^x[343]^x[335]^x[333]^x[324]^x[323]^x[322]^x[281]^x[280]^x[279]^x[278]^x[270]^x[269]^x[268]^x[267]^x[258]^x[256]^x[216]^x[214]^x[210]^x[208]^x[206]^x[204]^x[199]^x[197]^x[195]^x[183]^x[177]^x[172]^x[171]^x[166]^x[160]^x[108]^x[103]^x[102]^x[77]^x[76]^x[66]^x[56]^x[54]^x[46]^x[44]^x[40]^x[39]^x[38]^x[37]^x[35]^x[34]^x[33]^x[32]^x[23]^x[12]^x[11]^x[0];
	x_new[75]=x[343]^x[342]^x[334]^x[332]^x[323]^x[322]^x[321]^x[280]^x[279]^x[278]^x[269]^x[267]^x[256]^x[215]^x[214]^x[209]^x[208]^x[205]^x[198]^x[197]^x[194]^x[182]^x[176]^x[171]^x[165]^x[107]^x[102]^x[101]^x[76]^x[75]^x[65]^x[55]^x[54]^x[45]^x[39]^x[38]^x[37]^x[34]^x[33]^x[32]^x[22]^x[11];
	x_new[74]=x[342]^x[341]^x[333]^x[331]^x[322]^x[321]^x[320]^x[279]^x[278]^x[277]^x[268]^x[267]^x[266]^x[256]^x[214]^x[208]^x[204]^x[202]^x[197]^x[193]^x[181]^x[175]^x[170]^x[164]^x[106]^x[101]^x[100]^x[75]^x[74]^x[64]^x[54]^x[44]^x[42]^x[38]^x[37]^x[36]^x[33]^x[32]^x[21]^x[10];
	x_new[73]=x[351]^x[341]^x[340]^x[332]^x[321]^x[320]^x[287]^x[286]^x[278]^x[277]^x[275]^x[267]^x[265]^x[221]^x[213]^x[212]^x[211]^x[203]^x[199]^x[192]^x[180]^x[174]^x[169]^x[163]^x[122]^x[105]^x[99]^x[95]^x[73]^x[53]^x[52]^x[51]^x[47]^x[46]^x[45]^x[43]^x[41]^x[37]^x[35]^x[32]^x[20]^x[9];
	x_new[72]=x[351]^x[350]^x[340]^x[339]^x[331]^x[330]^x[320]^x[285]^x[277]^x[276]^x[275]^x[274]^x[266]^x[264]^x[223]^x[220]^x[212]^x[211]^x[210]^x[198]^x[179]^x[173]^x[168]^x[162]^x[104]^x[98]^x[94]^x[72]^x[63]^x[57]^x[52]^x[50]^x[46]^x[44]^x[40]^x[34]^x[19]^x[8];
	x_new[71]=x[373]^x[362]^x[351]^x[350]^x[349]^x[339]^x[338]^x[329]^x[284]^x[276]^x[275]^x[274]^x[273]^x[265]^x[263]^x[222]^x[219]^x[211]^x[210]^x[209]^x[197]^x[178]^x[172]^x[167]^x[161]^x[138]^x[132]^x[103]^x[97]^x[93]^x[71]^x[62]^x[56]^x[51]^x[49]^x[45]^x[43]^x[39]^x[33]^x[18]^x[7];
	x_new[70]=x[372]^x[361]^x[350]^x[349]^x[348]^x[338]^x[337]^x[328]^x[283]^x[275]^x[274]^x[273]^x[272]^x[264]^x[262]^x[221]^x[218]^x[210]^x[209]^x[208]^x[196]^x[177]^x[171]^x[166]^x[160]^x[137]^x[131]^x[102]^x[96]^x[92]^x[70]^x[61]^x[55]^x[50]^x[48]^x[44]^x[42]^x[38]^x[32]^x[17]^x[6];
	x_new[69]=x[371]^x[360]^x[349]^x[348]^x[347]^x[337]^x[336]^x[327]^x[282]^x[274]^x[273]^x[271]^x[263]^x[245]^x[234]^x[220]^x[217]^x[214]^x[209]^x[207]^x[197]^x[195]^x[192]^x[176]^x[165]^x[136]^x[130]^x[118]^x[108]^x[107]^x[106]^x[101]^x[97]^x[96]^x[91]^x[69]^x[60]^x[49]^x[47]^x[43]^x[41]^x[32]^x[16]^x[10]^x[5]^x[4];
	x_new[68]=x[370]^x[359]^x[348]^x[347]^x[346]^x[336]^x[335]^x[326]^x[281]^x[273]^x[272]^x[271]^x[270]^x[262]^x[260]^x[244]^x[233]^x[219]^x[216]^x[213]^x[208]^x[206]^x[202]^x[196]^x[194]^x[175]^x[164]^x[135]^x[129]^x[107]^x[106]^x[105]^x[100]^x[96]^x[90]^x[68]^x[59]^x[48]^x[46]^x[40]^x[36]^x[15]^x[9]^x[4]^x[3];
	x_new[67]=x[369]^x[358]^x[347]^x[346]^x[345]^x[335]^x[334]^x[325]^x[280]^x[272]^x[271]^x[270]^x[269]^x[261]^x[259]^x[243]^x[232]^x[218]^x[215]^x[212]^x[207]^x[205]^x[201]^x[195]^x[193]^x[174]^x[163]^x[134]^x[128]^x[106]^x[105]^x[104]^x[99]^x[89]^x[67]^x[58]^x[47]^x[45]^x[39]^x[35]^x[14]^x[8]^x[3]^x[2];
	x_new[66]=x[368]^x[357]^x[346]^x[345]^x[344]^x[334]^x[333]^x[324]^x[279]^x[271]^x[270]^x[269]^x[268]^x[260]^x[258]^x[242]^x[231]^x[217]^x[214]^x[211]^x[206]^x[204]^x[200]^x[194]^x[192]^x[173]^x[162]^x[133]^x[105]^x[104]^x[103]^x[98]^x[88]^x[66]^x[57]^x[46]^x[44]^x[38]^x[34]^x[13]^x[7]^x[2]^x[1];
	x_new[65]=x[345]^x[344]^x[343]^x[333]^x[332]^x[323]^x[278]^x[270]^x[269]^x[268]^x[267]^x[259]^x[257]^x[241]^x[230]^x[216]^x[210]^x[205]^x[203]^x[199]^x[193]^x[172]^x[161]^x[104]^x[103]^x[102]^x[97]^x[87]^x[65]^x[56]^x[45]^x[43]^x[37]^x[33]^x[12]^x[6]^x[1]^x[0];
	x_new[64]=x[344]^x[343]^x[342]^x[332]^x[331]^x[322]^x[278]^x[269]^x[268]^x[267]^x[258]^x[240]^x[229]^x[215]^x[209]^x[204]^x[203]^x[198]^x[171]^x[160]^x[103]^x[102]^x[101]^x[96]^x[86]^x[64]^x[55]^x[44]^x[43]^x[37]^x[11]^x[5]^x[0];
	x_new[63]=x[383]^x[373]^x[372]^x[371]^x[363]^x[361]^x[352]^x[333]^x[322]^x[311]^x[306]^x[301]^x[298]^x[295]^x[290]^x[288]^x[284]^x[278]^x[273]^x[267]^x[255]^x[254]^x[247]^x[246]^x[245]^x[244]^x[243]^x[235]^x[225]^x[186]^x[185]^x[181]^x[176]^x[174]^x[172]^x[171]^x[170]^x[167]^x[165]^x[161]^x[124]^x[113]^x[98]^x[95]^x[91]^x[90]^x[89]^x[80]^x[71]^x[70]^x[65]^x[63]^x[53]^x[49]^x[43]^x[37]^x[32]^x[26]^x[25]^x[21]^x[20]^x[19]^x[16]^x[15]^x[13]^x[12]^x[11]^x[6]^x[1]^x[0];
	x_new[62]=x[383]^x[382]^x[372]^x[371]^x[370]^x[360]^x[319]^x[310]^x[305]^x[300]^x[298]^x[297]^x[294]^x[289]^x[283]^x[277]^x[272]^x[266]^x[254]^x[253]^x[246]^x[245]^x[244]^x[242]^x[234]^x[233]^x[224]^x[190]^x[189]^x[178]^x[171]^x[170]^x[166]^x[160]^x[123]^x[112]^x[94]^x[88]^x[70]^x[69]^x[64]^x[63]^x[62]^x[52]^x[48]^x[36]^x[30]^x[24]^x[18]^x[12]^x[11]^x[10]^x[5]^x[4]^x[0];
	x_new[61]=x[382]^x[381]^x[371]^x[370]^x[369]^x[359]^x[342]^x[320]^x[318]^x[309]^x[304]^x[299]^x[297]^x[296]^x[293]^x[288]^x[282]^x[276]^x[271]^x[265]^x[255]^x[254]^x[253]^x[252]^x[245]^x[244]^x[241]^x[234]^x[233]^x[232]^x[191]^x[189]^x[188]^x[177]^x[169]^x[165]^x[122]^x[111]^x[107]^x[101]^x[96]^x[93]^x[87]^x[69]^x[62]^x[61]^x[51]^x[47]^x[35]^x[31]^x[29]^x[25]^x[23]^x[19]^x[17]^x[13]^x[11]^x[9]^x[3];
	x_new[60]=x[381]^x[380]^x[370]^x[369]^x[368]^x[358]^x[341]^x[330]^x[319]^x[317]^x[308]^x[303]^x[296]^x[295]^x[292]^x[281]^x[275]^x[270]^x[264]^x[254]^x[253]^x[252]^x[251]^x[244]^x[243]^x[240]^x[233]^x[232]^x[231]^x[190]^x[188]^x[187]^x[176]^x[168]^x[164]^x[121]^x[110]^x[106]^x[100]^x[92]^x[86]^x[68]^x[61]^x[60]^x[50]^x[46]^x[34]^x[30]^x[28]^x[24]^x[22]^x[18]^x[16]^x[12]^x[10]^x[8]^x[2];
	x_new[59]=x[380]^x[379]^x[369]^x[368]^x[367]^x[357]^x[340]^x[329]^x[318]^x[316]^x[307]^x[302]^x[295]^x[294]^x[291]^x[280]^x[274]^x[269]^x[263]^x[253]^x[252]^x[251]^x[250]^x[243]^x[242]^x[239]^x[232]^x[231]^x[230]^x[189]^x[187]^x[186]^x[175]^x[167]^x[163]^x[120]^x[109]^x[105]^x[99]^x[91]^x[85]^x[67]^x[60]^x[59]^x[49]^x[45]^x[33]^x[29]^x[27]^x[23]^x[21]^x[17]^x[15]^x[11]^x[9]^x[7]^x[1];
	x_new[58]=x[383]^x[379]^x[378]^x[377]^x[368]^x[367]^x[366]^x[356]^x[349]^x[339]^x[328]^x[317]^x[315]^x[306]^x[301]^x[294]^x[293]^x[290]^x[279]^x[273]^x[268]^x[262]^x[252]^x[251]^x[249]^x[242]^x[241]^x[238]^x[231]^x[230]^x[229]^x[223]^x[191]^x[190]^x[188]^x[184]^x[181]^x[180]^x[179]^x[175]^x[173]^x[171]^x[166]^x[162]^x[160]^x[147]^x[125]^x[108]^x[95]^x[90]^x[86]^x[85]^x[84]^x[75]^x[74]^x[66]^x[59]^x[58]^x[48]^x[44]^x[32]^x[31]^x[30]^x[28]^x[22]^x[21]^x[20]^x[19]^x[16]^x[14]^x[11]^x[10]^x[8]^x[6]^x[5];
	x_new[57]=x[382]^x[378]^x[377]^x[376]^x[367]^x[366]^x[365]^x[355]^x[348]^x[316]^x[314]^x[305]^x[300]^x[293]^x[292]^x[289]^x[278]^x[272]^x[267]^x[261]^x[251]^x[250]^x[249]^x[248]^x[241]^x[240]^x[237]^x[230]^x[229]^x[228]^x[222]^x[189]^x[187]^x[185]^x[184]^x[183]^x[180]^x[178]^x[174]^x[173]^x[172]^x[165]^x[161]^x[146]^x[124]^x[107]^x[103]^x[97]^x[95]^x[94]^x[89]^x[84]^x[83]^x[74]^x[73]^x[65]^x[58]^x[57]^x[47]^x[43]^x[29]^x[27]^x[25]^x[21]^x[20]^x[19]^x[18]^x[15]^x[13]^x[9]^x[7]^x[5];
	x_new[56]=x[381]^x[377]^x[376]^x[375]^x[366]^x[365]^x[364]^x[354]^x[347]^x[315]^x[313]^x[304]^x[299]^x[292]^x[291]^x[288]^x[277]^x[271]^x[266]^x[260]^x[250]^x[249]^x[248]^x[247]^x[240]^x[239]^x[236]^x[229]^x[228]^x[227]^x[221]^x[188]^x[186]^x[184]^x[183]^x[182]^x[179]^x[177]^x[173]^x[172]^x[171]^x[164]^x[160]^x[145]^x[123]^x[106]^x[102]^x[96]^x[95]^x[94]^x[93]^x[88]^x[83]^x[82]^x[74]^x[73]^x[72]^x[64]^x[57]^x[56]^x[46]^x[42]^x[28]^x[26]^x[24]^x[20]^x[19]^x[18]^x[17]^x[14]^x[12]^x[8]^x[6]^x[4];
	x_new[55]=x[380]^x[376]^x[375]^x[374]^x[365]^x[364]^x[363]^x[353]^x[346]^x[336]^x[325]^x[314]^x[312]^x[303]^x[291]^x[290]^x[276]^x[270]^x[265]^x[259]^x[249]^x[248]^x[247]^x[246]^x[239]^x[238]^x[235]^x[228]^x[227]^x[226]^x[220]^x[187]^x[185]^x[183]^x[181]^x[178]^x[176]^x[172]^x[170]^x[163]^x[144]^x[122]^x[105]^x[94]^x[93]^x[92]^x[87]^x[82]^x[81]^x[73]^x[72]^x[71]^x[56]^x[55]^x[45]^x[41]^x[27]^x[25]^x[23]^x[19]^x[18]^x[17]^x[16]^x[13]^x[11]^x[7]^x[5]^x[3];
	x_new[54]=x[379]^x[375]^x[374]^x[373]^x[364]^x[363]^x[362]^x[352]^x[345]^x[335]^x[324]^x[313]^x[311]^x[302]^x[290]^x[289]^x[275]^x[269]^x[264]^x[258]^x[248]^x[247]^x[246]^x[245]^x[238]^x[237]^x[234]^x[227]^x[226]^x[225]^x[219]^x[186]^x[184]^x[182]^x[180]^x[177]^x[175]^x[171]^x[169]^x[162]^x[143]^x[121]^x[104]^x[93]^x[92]^x[91]^x[86]^x[81]^x[80]^x[72]^x[71]^x[70]^x[55]^x[54]^x[44]^x[40]^x[26]^x[24]^x[22]^x[18]^x[17]^x[16]^x[15]^x[12]^x[10]^x[6]^x[4]^x[2];
	x_new[53]=x[378]^x[374]^x[373]^x[372]^x[363]^x[361]^x[344]^x[334]^x[323]^x[312]^x[310]^x[301]^x[289]^x[288]^x[274]^x[268]^x[263]^x[257]^x[247]^x[244]^x[237]^x[236]^x[234]^x[233]^x[226]^x[225]^x[218]^x[185]^x[183]^x[181]^x[179]^x[176]^x[174]^x[171]^x[168]^x[161]^x[160]^x[142]^x[120]^x[103]^x[92]^x[91]^x[90]^x[85]^x[80]^x[79]^x[71]^x[70]^x[69]^x[54]^x[53]^x[43]^x[39]^x[25]^x[23]^x[21]^x[17]^x[16]^x[15]^x[14]^x[10]^x[9]^x[4]^x[3]^x[1]^x[0];
	x_new[52]=x[382]^x[373]^x[372]^x[362]^x[360]^x[333]^x[322]^x[319]^x[311]^x[309]^x[300]^x[298]^x[288]^x[273]^x[267]^x[262]^x[256]^x[255]^x[254]^x[246]^x[243]^x[236]^x[235]^x[232]^x[225]^x[224]^x[191]^x[190]^x[186]^x[185]^x[182]^x[180]^x[178]^x[174]^x[169]^x[160]^x[113]^x[102]^x[98]^x[91]^x[90]^x[84]^x[80]^x[78]^x[70]^x[53]^x[52]^x[42]^x[38]^x[31]^x[30]^x[26]^x[24]^x[22]^x[16]^x[14]^x[10]^x[9]^x[8]^x[4]^x[3]^x[2]^x[0];
	x_new[51]=x[381]^x[372]^x[371]^x[361]^x[359]^x[319]^x[318]^x[310]^x[308]^x[299]^x[298]^x[297]^x[272]^x[261]^x[255]^x[254]^x[253]^x[245]^x[244]^x[243]^x[242]^x[235]^x[233]^x[231]^x[224]^x[191]^x[189]^x[181]^x[178]^x[177]^x[170]^x[168]^x[167]^x[112]^x[101]^x[90]^x[83]^x[77]^x[69]^x[52]^x[51]^x[41]^x[37]^x[31]^x[29]^x[25]^x[23]^x[21]^x[19]^x[15]^x[13]^x[10]^x[9]^x[8]^x[7]^x[4]^x[3]^x[2]^x[1];
	x_new[50]=x[380]^x[371]^x[370]^x[360]^x[358]^x[318]^x[317]^x[309]^x[307]^x[298]^x[297]^x[296]^x[271]^x[260]^x[255]^x[254]^x[253]^x[252]^x[244]^x[243]^x[242]^x[241]^x[232]^x[230]^x[190]^x[188]^x[180]^x[177]^x[176]^x[169]^x[167]^x[166]^x[111]^x[100]^x[82]^x[76]^x[51]^x[50]^x[40]^x[36]^x[30]^x[28]^x[24]^x[22]^x[20]^x[18]^x[14]^x[12]^x[9]^x[8]^x[7]^x[6]^x[3]^x[2]^x[1]^x[0];
	x_new[49]=x[379]^x[370]^x[369]^x[359]^x[357]^x[317]^x[316]^x[308]^x[306]^x[297]^x[296]^x[295]^x[270]^x[259]^x[254]^x[253]^x[252]^x[251]^x[243]^x[242]^x[241]^x[240]^x[231]^x[229]^x[189]^x[187]^x[182]^x[181]^x[179]^x[170]^x[168]^x[166]^x[164]^x[160]^x[138]^x[110]^x[99]^x[81]^x[75]^x[50]^x[49]^x[39]^x[35]^x[29]^x[27]^x[23]^x[22]^x[19]^x[17]^x[13]^x[11]^x[10]^x[8]^x[7]^x[6]^x[5]^x[2]^x[1];
	x_new[48]=x[378]^x[369]^x[368]^x[358]^x[356]^x[316]^x[315]^x[307]^x[305]^x[296]^x[295]^x[294]^x[269]^x[258]^x[253]^x[252]^x[251]^x[250]^x[242]^x[241]^x[240]^x[239]^x[230]^x[228]^x[188]^x[186]^x[180]^x[178]^x[175]^x[169]^x[167]^x[165]^x[164]^x[163]^x[137]^x[109]^x[98]^x[80]^x[74]^x[49]^x[48]^x[38]^x[34]^x[28]^x[26]^x[22]^x[18]^x[16]^x[12]^x[10]^x[9]^x[7]^x[6]^x[5]^x[4]^x[1]^x[0];
	x_new[47]=x[377]^x[368]^x[367]^x[357]^x[355]^x[315]^x[314]^x[306]^x[304]^x[295]^x[294]^x[293]^x[268]^x[257]^x[252]^x[251]^x[250]^x[249]^x[241]^x[240]^x[239]^x[238]^x[229]^x[227]^x[187]^x[185]^x[181]^x[179]^x[177]^x[175]^x[174]^x[170]^x[168]^x[166]^x[163]^x[162]^x[136]^x[108]^x[97]^x[79]^x[75]^x[74]^x[73]^x[64]^x[48]^x[47]^x[37]^x[33]^x[27]^x[25]^x[17]^x[15]^x[11]^x[10]^x[9]^x[8]^x[6]^x[5]^x[4]^x[3]^x[0];
	x_new[46]=x[376]^x[367]^x[366]^x[356]^x[354]^x[314]^x[313]^x[305]^x[303]^x[294]^x[293]^x[292]^x[267]^x[256]^x[251]^x[250]^x[249]^x[248]^x[240]^x[239]^x[238]^x[237]^x[228]^x[226]^x[186]^x[184]^x[180]^x[178]^x[176]^x[174]^x[173]^x[169]^x[167]^x[165]^x[162]^x[161]^x[135]^x[107]^x[96]^x[78]^x[73]^x[72]^x[47]^x[46]^x[36]^x[32]^x[26]^x[24]^x[16]^x[14]^x[10]^x[9]^x[8]^x[7]^x[5]^x[4]^x[3]^x[2];
	x_new[45]=x[375]^x[366]^x[365]^x[355]^x[353]^x[313]^x[312]^x[304]^x[302]^x[293]^x[292]^x[291]^x[250]^x[249]^x[248]^x[247]^x[239]^x[238]^x[237]^x[236]^x[227]^x[225]^x[185]^x[183]^x[179]^x[177]^x[175]^x[173]^x[172]^x[168]^x[166]^x[164]^x[161]^x[160]^x[134]^x[77]^x[72]^x[71]^x[46]^x[45]^x[35]^x[25]^x[23]^x[15]^x[13]^x[9]^x[8]^x[7]^x[6]^x[4]^x[3]^x[2]^x[1];
	x_new[44]=x[374]^x[365]^x[364]^x[354]^x[352]^x[312]^x[311]^x[303]^x[301]^x[292]^x[291]^x[290]^x[249]^x[248]^x[247]^x[246]^x[238]^x[237]^x[236]^x[235]^x[226]^x[224]^x[184]^x[182]^x[178]^x[176]^x[174]^x[172]^x[167]^x[165]^x[163]^x[133]^x[76]^x[71]^x[70]^x[45]^x[44]^x[34]^x[24]^x[22]^x[14]^x[12]^x[8]^x[7]^x[6]^x[5]^x[3]^x[2]^x[1]^x[0];
	x_new[43]=x[364]^x[363]^x[353]^x[311]^x[310]^x[302]^x[300]^x[291]^x[290]^x[289]^x[248]^x[247]^x[246]^x[237]^x[235]^x[224]^x[183]^x[182]^x[177]^x[176]^x[173]^x[166]^x[165]^x[162]^x[75]^x[70]^x[69]^x[44]^x[43]^x[33]^x[23]^x[22]^x[13]^x[7]^x[6]^x[5]^x[2]^x[1]^x[0];
	x_new[42]=x[363]^x[362]^x[352]^x[310]^x[309]^x[301]^x[299]^x[290]^x[289]^x[288]^x[247]^x[246]^x[245]^x[236]^x[235]^x[234]^x[224]^x[182]^x[176]^x[172]^x[170]^x[165]^x[161]^x[74]^x[69]^x[68]^x[43]^x[42]^x[32]^x[22]^x[12]^x[10]^x[6]^x[5]^x[4]^x[1]^x[0];
	x_new[41]=x[383]^x[361]^x[319]^x[309]^x[308]^x[300]^x[289]^x[288]^x[255]^x[254]^x[246]^x[245]^x[243]^x[235]^x[233]^x[189]^x[181]^x[180]^x[179]^x[171]^x[167]^x[160]^x[90]^x[73]^x[67]^x[63]^x[41]^x[21]^x[20]^x[19]^x[15]^x[14]^x[13]^x[11]^x[9]^x[5]^x[3]^x[0];
	x_new[40]=x[382]^x[360]^x[319]^x[318]^x[308]^x[307]^x[299]^x[298]^x[288]^x[253]^x[245]^x[244]^x[243]^x[242]^x[234]^x[232]^x[191]^x[188]^x[180]^x[179]^x[178]^x[166]^x[72]^x[66]^x[62]^x[40]^x[31]^x[25]^x[20]^x[18]^x[14]^x[12]^x[8]^x[2];
	x_new[39]=x[381]^x[359]^x[341]^x[330]^x[319]^x[318]^x[317]^x[307]^x[306]^x[297]^x[252]^x[244]^x[243]^x[242]^x[241]^x[233]^x[231]^x[190]^x[187]^x[179]^x[178]^x[177]^x[165]^x[106]^x[100]^x[71]^x[65]^x[61]^x[39]^x[30]^x[24]^x[19]^x[17]^x[13]^x[11]^x[7]^x[1];
	x_new[38]=x[380]^x[358]^x[340]^x[329]^x[318]^x[317]^x[316]^x[306]^x[305]^x[296]^x[251]^x[243]^x[242]^x[241]^x[240]^x[232]^x[230]^x[189]^x[186]^x[178]^x[177]^x[176]^x[164]^x[105]^x[99]^x[70]^x[64]^x[60]^x[38]^x[29]^x[23]^x[18]^x[16]^x[12]^x[10]^x[6]^x[0];
	x_new[37]=x[379]^x[373]^x[367]^x[362]^x[357]^x[356]^x[339]^x[328]^x[317]^x[316]^x[315]^x[305]^x[304]^x[295]^x[250]^x[242]^x[241]^x[239]^x[231]^x[213]^x[202]^x[188]^x[185]^x[182]^x[177]^x[175]^x[165]^x[163]^x[160]^x[104]^x[98]^x[86]^x[76]^x[75]^x[74]^x[69]^x[65]^x[64]^x[59]^x[37]^x[28]^x[17]^x[15]^x[11]^x[9]^x[0];
	x_new[36]=x[378]^x[372]^x[366]^x[361]^x[356]^x[355]^x[338]^x[327]^x[316]^x[315]^x[314]^x[304]^x[303]^x[294]^x[249]^x[241]^x[240]^x[239]^x[238]^x[230]^x[228]^x[212]^x[201]^x[187]^x[184]^x[181]^x[176]^x[174]^x[170]^x[164]^x[162]^x[103]^x[97]^x[75]^x[74]^x[73]^x[68]^x[64]^x[58]^x[36]^x[27]^x[16]^x[14]^x[8]^x[4];
	x_new[35]=x[377]^x[371]^x[365]^x[360]^x[355]^x[354]^x[337]^x[326]^x[315]^x[314]^x[313]^x[303]^x[302]^x[293]^x[248]^x[240]^x[239]^x[238]^x[237]^x[229]^x[227]^x[211]^x[200]^x[186]^x[183]^x[180]^x[175]^x[173]^x[169]^x[163]^x[161]^x[102]^x[96]^x[74]^x[73]^x[72]^x[67]^x[57]^x[35]^x[26]^x[15]^x[13]^x[7]^x[3];
	x_new[34]=x[376]^x[370]^x[364]^x[359]^x[354]^x[353]^x[336]^x[325]^x[314]^x[313]^x[312]^x[302]^x[301]^x[292]^x[247]^x[239]^x[238]^x[237]^x[236]^x[228]^x[226]^x[210]^x[199]^x[185]^x[182]^x[179]^x[174]^x[172]^x[168]^x[162]^x[160]^x[101]^x[73]^x[72]^x[71]^x[66]^x[56]^x[34]^x[25]^x[14]^x[12]^x[6]^x[2];
	x_new[33]=x[375]^x[369]^x[363]^x[358]^x[353]^x[352]^x[313]^x[312]^x[311]^x[301]^x[300]^x[291]^x[246]^x[238]^x[237]^x[236]^x[235]^x[227]^x[225]^x[209]^x[198]^x[184]^x[178]^x[173]^x[171]^x[167]^x[161]^x[72]^x[71]^x[70]^x[65]^x[55]^x[33]^x[24]^x[13]^x[11]^x[5]^x[1];
	x_new[32]=x[374]^x[368]^x[357]^x[352]^x[312]^x[311]^x[310]^x[300]^x[299]^x[290]^x[246]^x[237]^x[236]^x[235]^x[226]^x[208]^x[197]^x[183]^x[177]^x[172]^x[171]^x[166]^x[71]^x[70]^x[69]^x[64]^x[54]^x[32]^x[23]^x[12]^x[11]^x[5];
	x_new[31]=x[383]^x[382]^x[379]^x[377]^x[376]^x[375]^x[374]^x[373]^x[372]^x[371]^x[369]^x[365]^x[363]^x[358]^x[357]^x[356]^x[353]^x[351]^x[341]^x[340]^x[339]^x[331]^x[329]^x[320]^x[301]^x[290]^x[279]^x[274]^x[269]^x[266]^x[263]^x[258]^x[256]^x[252]^x[246]^x[241]^x[235]^x[223]^x[222]^x[215]^x[214]^x[213]^x[212]^x[211]^x[203]^x[193]^x[137]^x[92]^x[81]^x[66]^x[63]^x[59]^x[58]^x[57]^x[48]^x[39]^x[38]^x[33]^x[31]^x[21]^x[17]^x[11]^x[5]^x[0];
	x_new[30]=x[382]^x[381]^x[376]^x[375]^x[374]^x[373]^x[372]^x[370]^x[368]^x[367]^x[366]^x[364]^x[362]^x[361]^x[357]^x[356]^x[355]^x[352]^x[351]^x[350]^x[340]^x[339]^x[338]^x[328]^x[287]^x[278]^x[273]^x[268]^x[266]^x[265]^x[262]^x[257]^x[251]^x[245]^x[240]^x[234]^x[222]^x[221]^x[214]^x[213]^x[212]^x[210]^x[202]^x[201]^x[192]^x[157]^x[146]^x[91]^x[80]^x[62]^x[56]^x[38]^x[37]^x[32]^x[31]^x[30]^x[20]^x[16]^x[4];
	x_new[29]=x[383]^x[382]^x[381]^x[380]^x[377]^x[376]^x[375]^x[374]^x[373]^x[372]^x[369]^x[367]^x[366]^x[363]^x[362]^x[361]^x[360]^x[356]^x[355]^x[354]^x[350]^x[349]^x[339]^x[338]^x[337]^x[327]^x[310]^x[288]^x[286]^x[277]^x[272]^x[267]^x[265]^x[264]^x[261]^x[256]^x[250]^x[244]^x[239]^x[233]^x[223]^x[222]^x[221]^x[220]^x[213]^x[212]^x[209]^x[202]^x[201]^x[200]^x[156]^x[145]^x[135]^x[90]^x[79]^x[75]^x[69]^x[64]^x[61]^x[55]^x[37]^x[30]^x[29]^x[19]^x[15]^x[3];
	x_new[28]=x[382]^x[381]^x[380]^x[379]^x[376]^x[375]^x[374]^x[373]^x[372]^x[371]^x[368]^x[366]^x[365]^x[362]^x[361]^x[360]^x[359]^x[355]^x[354]^x[353]^x[349]^x[348]^x[338]^x[337]^x[336]^x[326]^x[309]^x[298]^x[287]^x[285]^x[276]^x[271]^x[264]^x[263]^x[260]^x[249]^x[243]^x[238]^x[232]^x[222]^x[221]^x[220]^x[219]^x[212]^x[211]^x[208]^x[201]^x[200]^x[199]^x[155]^x[144]^x[134]^x[89]^x[78]^x[74]^x[68]^x[60]^x[54]^x[36]^x[29]^x[28]^x[18]^x[14]^x[2];
	x_new[27]=x[381]^x[380]^x[379]^x[378]^x[375]^x[374]^x[373]^x[372]^x[371]^x[370]^x[367]^x[365]^x[364]^x[361]^x[360]^x[359]^x[358]^x[354]^x[353]^x[352]^x[348]^x[347]^x[337]^x[336]^x[335]^x[325]^x[308]^x[297]^x[286]^x[284]^x[275]^x[270]^x[263]^x[262]^x[259]^x[248]^x[242]^x[237]^x[231]^x[221]^x[220]^x[219]^x[218]^x[211]^x[210]^x[207]^x[200]^x[199]^x[198]^x[154]^x[143]^x[133]^x[88]^x[77]^x[73]^x[67]^x[59]^x[53]^x[35]^x[28]^x[27]^x[17]^x[13]^x[1];
	x_new[26]=x[380]^x[379]^x[377]^x[373]^x[370]^x[369]^x[366]^x[364]^x[361]^x[360]^x[359]^x[358]^x[357]^x[353]^x[352]^x[351]^x[347]^x[346]^x[345]^x[336]^x[335]^x[334]^x[324]^x[317]^x[307]^x[296]^x[285]^x[283]^x[274]^x[269]^x[262]^x[261]^x[258]^x[247]^x[241]^x[236]^x[230]^x[220]^x[219]^x[217]^x[210]^x[209]^x[206]^x[199]^x[198]^x[197]^x[191]^x[153]^x[132]^x[115]^x[93]^x[76]^x[63]^x[58]^x[54]^x[53]^x[52]^x[43]^x[42]^x[34]^x[27]^x[26]^x[16]^x[12]^x[0];
	x_new[25]=x[383]^x[382]^x[379]^x[378]^x[377]^x[376]^x[373]^x[369]^x[368]^x[365]^x[363]^x[361]^x[360]^x[359]^x[358]^x[357]^x[356]^x[352]^x[350]^x[346]^x[345]^x[344]^x[335]^x[334]^x[333]^x[323]^x[316]^x[284]^x[282]^x[273]^x[268]^x[261]^x[260]^x[257]^x[246]^x[240]^x[235]^x[229]^x[219]^x[218]^x[217]^x[216]^x[209]^x[208]^x[205]^x[198]^x[197]^x[196]^x[190]^x[152]^x[141]^x[131]^x[114]^x[92]^x[75]^x[71]^x[65]^x[63]^x[62]^x[57]^x[52]^x[51]^x[42]^x[41]^x[33]^x[26]^x[25]^x[15]^x[11];
	x_new[24]=x[383]^x[382]^x[381]^x[378]^x[377]^x[376]^x[375]^x[372]^x[368]^x[367]^x[364]^x[360]^x[359]^x[358]^x[357]^x[356]^x[355]^x[349]^x[345]^x[344]^x[343]^x[334]^x[333]^x[332]^x[322]^x[315]^x[283]^x[281]^x[272]^x[267]^x[260]^x[259]^x[256]^x[245]^x[239]^x[234]^x[228]^x[218]^x[217]^x[216]^x[215]^x[208]^x[207]^x[204]^x[197]^x[196]^x[195]^x[189]^x[151]^x[140]^x[130]^x[113]^x[91]^x[74]^x[70]^x[64]^x[63]^x[62]^x[61]^x[56]^x[51]^x[50]^x[42]^x[41]^x[40]^x[32]^x[25]^x[24]^x[14]^x[10];
	x_new[23]=x[382]^x[381]^x[380]^x[377]^x[376]^x[375]^x[374]^x[371]^x[367]^x[366]^x[363]^x[359]^x[358]^x[357]^x[356]^x[355]^x[354]^x[348]^x[344]^x[343]^x[342]^x[333]^x[332]^x[331]^x[321]^x[314]^x[304]^x[293]^x[282]^x[280]^x[271]^x[259]^x[258]^x[244]^x[238]^x[233]^x[227]^x[217]^x[216]^x[215]^x[214]^x[207]^x[206]^x[203]^x[196]^x[195]^x[194]^x[188]^x[129]^x[112]^x[90]^x[73]^x[62]^x[61]^x[60]^x[55]^x[50]^x[49]^x[41]^x[40]^x[39]^x[24]^x[23]^x[13]^x[9];
	x_new[22]=x[381]^x[380]^x[379]^x[376]^x[375]^x[374]^x[373]^x[370]^x[366]^x[365]^x[362]^x[358]^x[357]^x[356]^x[355]^x[354]^x[353]^x[347]^x[343]^x[342]^x[341]^x[332]^x[331]^x[330]^x[320]^x[313]^x[303]^x[292]^x[281]^x[279]^x[270]^x[258]^x[257]^x[243]^x[237]^x[232]^x[226]^x[216]^x[215]^x[214]^x[213]^x[206]^x[205]^x[202]^x[195]^x[194]^x[193]^x[187]^x[128]^x[111]^x[89]^x[72]^x[61]^x[60]^x[59]^x[54]^x[49]^x[48]^x[40]^x[39]^x[38]^x[23]^x[22]^x[12]^x[8];
	x_new[21]=x[380]^x[379]^x[378]^x[375]^x[372]^x[369]^x[368]^x[367]^x[365]^x[364]^x[362]^x[361]^x[355]^x[354]^x[353]^x[346]^x[342]^x[341]^x[340]^x[331]^x[329]^x[312]^x[302]^x[291]^x[280]^x[278]^x[269]^x[257]^x[256]^x[242]^x[236]^x[231]^x[225]^x[215]^x[212]^x[205]^x[204]^x[202]^x[201]^x[194]^x[193]^x[186]^x[110]^x[88]^x[71]^x[60]^x[59]^x[58]^x[53]^x[48]^x[47]^x[39]^x[38]^x[37]^x[22]^x[21]^x[11]^x[7];
	x_new[20]=x[383]^x[382]^x[379]^x[378]^x[377]^x[376]^x[374]^x[371]^x[367]^x[366]^x[365]^x[364]^x[363]^x[360]^x[357]^x[356]^x[354]^x[353]^x[352]^x[350]^x[341]^x[340]^x[330]^x[328]^x[301]^x[290]^x[287]^x[279]^x[277]^x[268]^x[266]^x[256]^x[241]^x[235]^x[230]^x[224]^x[223]^x[222]^x[214]^x[211]^x[204]^x[203]^x[200]^x[193]^x[192]^x[81]^x[70]^x[66]^x[59]^x[58]^x[52]^x[48]^x[46]^x[38]^x[21]^x[20]^x[10]^x[6];
	x_new[19]=x[383]^x[382]^x[381]^x[378]^x[377]^x[376]^x[375]^x[373]^x[372]^x[371]^x[370]^x[367]^x[366]^x[365]^x[364]^x[363]^x[361]^x[359]^x[355]^x[353]^x[352]^x[349]^x[340]^x[339]^x[329]^x[327]^x[287]^x[286]^x[278]^x[276]^x[267]^x[266]^x[265]^x[240]^x[229]^x[223]^x[222]^x[221]^x[213]^x[212]^x[211]^x[210]^x[203]^x[201]^x[199]^x[192]^x[146]^x[135]^x[80]^x[69]^x[58]^x[51]^x[45]^x[37]^x[20]^x[19]^x[9]^x[5];
	x_new[18]=x[383]^x[382]^x[381]^x[380]^x[377]^x[376]^x[375]^x[374]^x[372]^x[371]^x[370]^x[369]^x[366]^x[365]^x[364]^x[363]^x[360]^x[358]^x[354]^x[352]^x[348]^x[339]^x[338]^x[328]^x[326]^x[286]^x[285]^x[277]^x[275]^x[266]^x[265]^x[264]^x[239]^x[228]^x[223]^x[222]^x[221]^x[220]^x[212]^x[211]^x[210]^x[209]^x[200]^x[198]^x[145]^x[134]^x[79]^x[68]^x[50]^x[44]^x[19]^x[18]^x[8]^x[4];
	x_new[17]=x[382]^x[381]^x[380]^x[379]^x[376]^x[375]^x[373]^x[371]^x[370]^x[369]^x[368]^x[365]^x[363]^x[362]^x[359]^x[357]^x[347]^x[338]^x[337]^x[327]^x[325]^x[285]^x[284]^x[276]^x[274]^x[265]^x[264]^x[263]^x[238]^x[227]^x[222]^x[221]^x[220]^x[219]^x[211]^x[210]^x[209]^x[208]^x[199]^x[197]^x[144]^x[106]^x[78]^x[67]^x[49]^x[43]^x[18]^x[17]^x[7]^x[3];
	x_new[16]=x[381]^x[380]^x[379]^x[378]^x[375]^x[374]^x[373]^x[372]^x[370]^x[369]^x[368]^x[367]^x[364]^x[363]^x[362]^x[361]^x[358]^x[356]^x[352]^x[346]^x[337]^x[336]^x[326]^x[324]^x[284]^x[283]^x[275]^x[273]^x[264]^x[263]^x[262]^x[237]^x[226]^x[221]^x[220]^x[219]^x[218]^x[210]^x[209]^x[208]^x[207]^x[198]^x[196]^x[143]^x[132]^x[105]^x[77]^x[66]^x[48]^x[42]^x[17]^x[16]^x[6]^x[2];
	x_new[15]=x[380]^x[379]^x[378]^x[377]^x[374]^x[373]^x[372]^x[371]^x[369]^x[368]^x[367]^x[366]^x[362]^x[361]^x[360]^x[357]^x[355]^x[352]^x[345]^x[336]^x[335]^x[325]^x[323]^x[283]^x[282]^x[274]^x[272]^x[263]^x[262]^x[261]^x[236]^x[225]^x[220]^x[219]^x[218]^x[217]^x[209]^x[208]^x[207]^x[206]^x[197]^x[195]^x[142]^x[131]^x[104]^x[76]^x[65]^x[47]^x[43]^x[42]^x[41]^x[32]^x[16]^x[15]^x[5]^x[1];
	x_new[14]=x[379]^x[378]^x[377]^x[376]^x[373]^x[372]^x[371]^x[370]^x[368]^x[367]^x[366]^x[365]^x[362]^x[361]^x[360]^x[359]^x[356]^x[354]^x[344]^x[335]^x[334]^x[324]^x[322]^x[282]^x[281]^x[273]^x[271]^x[262]^x[261]^x[260]^x[235]^x[224]^x[219]^x[218]^x[217]^x[216]^x[208]^x[207]^x[206]^x[205]^x[196]^x[194]^x[141]^x[130]^x[103]^x[75]^x[64]^x[46]^x[41]^x[40]^x[15]^x[14]^x[4]^x[0];
	x_new[13]=x[378]^x[377]^x[376]^x[375]^x[372]^x[371]^x[370]^x[369]^x[367]^x[366]^x[365]^x[364]^x[361]^x[360]^x[359]^x[358]^x[355]^x[353]^x[343]^x[334]^x[333]^x[323]^x[321]^x[281]^x[280]^x[272]^x[270]^x[261]^x[260]^x[259]^x[218]^x[217]^x[216]^x[215]^x[207]^x[206]^x[205]^x[204]^x[195]^x[193]^x[140]^x[129]^x[102]^x[45]^x[40]^x[39]^x[14]^x[13]^x[3];
	x_new[12]=x[377]^x[376]^x[375]^x[374]^x[371]^x[370]^x[369]^x[368]^x[366]^x[365]^x[364]^x[363]^x[360]^x[359]^x[358]^x[357]^x[354]^x[352]^x[342]^x[333]^x[332]^x[322]^x[320]^x[280]^x[279]^x[271]^x[269]^x[260]^x[259]^x[258]^x[217]^x[216]^x[215]^x[214]^x[206]^x[205]^x[204]^x[203]^x[194]^x[192]^x[101]^x[44]^x[39]^x[38]^x[13]^x[12]^x[2];
	x_new[11]=x[376]^x[375]^x[374]^x[370]^x[369]^x[368]^x[365]^x[363]^x[359]^x[358]^x[357]^x[352]^x[332]^x[331]^x[321]^x[279]^x[278]^x[270]^x[268]^x[259]^x[258]^x[257]^x[216]^x[215]^x[214]^x[205]^x[203]^x[192]^x[43]^x[38]^x[37]^x[12]^x[11]^x[1];
	x_new[10]=x[375]^x[374]^x[373]^x[369]^x[368]^x[367]^x[364]^x[363]^x[362]^x[358]^x[357]^x[356]^x[352]^x[331]^x[330]^x[320]^x[278]^x[277]^x[269]^x[267]^x[258]^x[257]^x[256]^x[215]^x[214]^x[213]^x[204]^x[203]^x[202]^x[192]^x[42]^x[37]^x[36]^x[11]^x[10]^x[0];
	x_new[9]=x[383]^x[382]^x[378]^x[377]^x[376]^x[374]^x[373]^x[371]^x[368]^x[367]^x[365]^x[363]^x[361]^x[357]^x[355]^x[351]^x[329]^x[287]^x[277]^x[276]^x[268]^x[257]^x[256]^x[223]^x[222]^x[214]^x[213]^x[211]^x[203]^x[201]^x[157]^x[136]^x[58]^x[41]^x[35]^x[31]^x[9];
	x_new[8]=x[381]^x[375]^x[373]^x[372]^x[371]^x[370]^x[367]^x[366]^x[365]^x[364]^x[362]^x[360]^x[356]^x[354]^x[350]^x[328]^x[287]^x[286]^x[276]^x[275]^x[267]^x[266]^x[256]^x[221]^x[213]^x[212]^x[211]^x[210]^x[202]^x[200]^x[156]^x[40]^x[34]^x[30]^x[8];
	x_new[7]=x[380]^x[374]^x[372]^x[371]^x[370]^x[369]^x[366]^x[365]^x[364]^x[363]^x[361]^x[359]^x[355]^x[353]^x[349]^x[327]^x[309]^x[298]^x[287]^x[286]^x[285]^x[275]^x[274]^x[265]^x[220]^x[212]^x[211]^x[210]^x[209]^x[201]^x[199]^x[155]^x[74]^x[68]^x[39]^x[33]^x[29]^x[7];
	x_new[6]=x[379]^x[373]^x[371]^x[370]^x[369]^x[368]^x[365]^x[364]^x[363]^x[362]^x[360]^x[358]^x[354]^x[352]^x[348]^x[326]^x[308]^x[297]^x[286]^x[285]^x[284]^x[274]^x[273]^x[264]^x[219]^x[211]^x[210]^x[209]^x[208]^x[200]^x[198]^x[154]^x[73]^x[67]^x[38]^x[32]^x[28]^x[6];
	x_new[5]=x[378]^x[374]^x[372]^x[370]^x[369]^x[367]^x[361]^x[359]^x[352]^x[347]^x[341]^x[335]^x[330]^x[325]^x[324]^x[307]^x[296]^x[285]^x[284]^x[283]^x[273]^x[272]^x[263]^x[218]^x[210]^x[209]^x[207]^x[199]^x[181]^x[170]^x[153]^x[72]^x[66]^x[54]^x[44]^x[43]^x[42]^x[37]^x[33]^x[32]^x[27]^x[5];
	x_new[4]=x[377]^x[371]^x[369]^x[368]^x[367]^x[366]^x[360]^x[358]^x[356]^x[346]^x[340]^x[334]^x[329]^x[324]^x[323]^x[306]^x[295]^x[284]^x[283]^x[282]^x[272]^x[271]^x[262]^x[217]^x[209]^x[208]^x[207]^x[206]^x[198]^x[196]^x[180]^x[169]^x[152]^x[71]^x[65]^x[43]^x[42]^x[41]^x[36]^x[32]^x[26]^x[4];
	x_new[3]=x[376]^x[370]^x[368]^x[367]^x[366]^x[365]^x[359]^x[357]^x[355]^x[345]^x[339]^x[333]^x[328]^x[323]^x[322]^x[305]^x[294]^x[283]^x[282]^x[281]^x[271]^x[270]^x[261]^x[216]^x[208]^x[207]^x[206]^x[205]^x[197]^x[195]^x[179]^x[168]^x[151]^x[70]^x[64]^x[42]^x[41]^x[40]^x[35]^x[25]^x[3];
	x_new[2]=x[375]^x[369]^x[367]^x[366]^x[365]^x[364]^x[358]^x[356]^x[354]^x[344]^x[338]^x[332]^x[327]^x[322]^x[321]^x[304]^x[293]^x[282]^x[281]^x[280]^x[270]^x[269]^x[260]^x[215]^x[207]^x[206]^x[205]^x[204]^x[196]^x[194]^x[178]^x[167]^x[150]^x[69]^x[41]^x[40]^x[39]^x[34]^x[24]^x[2];
	x_new[1]=x[374]^x[368]^x[366]^x[365]^x[364]^x[363]^x[357]^x[355]^x[353]^x[343]^x[337]^x[331]^x[326]^x[321]^x[320]^x[281]^x[280]^x[279]^x[269]^x[268]^x[259]^x[214]^x[206]^x[205]^x[204]^x[203]^x[195]^x[193]^x[177]^x[166]^x[40]^x[39]^x[38]^x[33]^x[23]^x[1];
	x_new[0]=x[374]^x[368]^x[365]^x[364]^x[363]^x[357]^x[354]^x[342]^x[336]^x[325]^x[320]^x[280]^x[279]^x[278]^x[268]^x[267]^x[258]^x[214]^x[205]^x[204]^x[203]^x[194]^x[176]^x[165]^x[39]^x[38]^x[37]^x[32]^x[22]^x[0];
	return x_new;
endfunction
endpackage
