function Bit#(330) encode(Bit#(330) x, Bit#(32) u);
	Bit#(330) y;
	y[0] = x[298]^x[299]^x[300]^x[301]^x[302]^x[304]^x[306]^x[307]^x[310]^x[316]^x[318]^x[319]^x[320]^x[323]^x[324]^x[325]^x[326]^x[327]^u[31]^u[30]^u[29]^u[28]^u[27]^u[25]^u[23]^u[22]^u[19]^u[13]^u[11]^u[10]^u[9]^u[6]^u[5]^u[4]^u[3]^u[2];
	y[1] = x[298]^x[303]^x[304]^x[305]^x[306]^x[308]^x[310]^x[311]^x[316]^x[317]^x[318]^x[321]^x[323]^x[328]^u[31]^u[26]^u[25]^u[24]^u[23]^u[21]^u[19]^u[18]^u[13]^u[12]^u[11]^u[8]^u[6]^u[1];
	y[2] = x[298]^x[300]^x[301]^x[302]^x[305]^x[309]^x[310]^x[311]^x[312]^x[316]^x[317]^x[320]^x[322]^x[323]^x[325]^x[326]^x[327]^x[329]^u[31]^u[29]^u[28]^u[27]^u[24]^u[20]^u[19]^u[18]^u[17]^u[13]^u[12]^u[9]^u[7]^u[6]^u[4]^u[3]^u[2]^u[0];
	y[3] = x[299]^x[301]^x[302]^x[303]^x[306]^x[310]^x[311]^x[312]^x[313]^x[317]^x[318]^x[321]^x[323]^x[324]^x[326]^x[327]^x[328]^u[30]^u[28]^u[27]^u[26]^u[23]^u[19]^u[18]^u[17]^u[16]^u[12]^u[11]^u[8]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[4] = x[298]^x[299]^x[301]^x[303]^x[306]^x[310]^x[311]^x[312]^x[313]^x[314]^x[316]^x[320]^x[322]^x[323]^x[326]^x[328]^x[329]^u[31]^u[30]^u[28]^u[26]^u[23]^u[19]^u[18]^u[17]^u[16]^u[15]^u[13]^u[9]^u[7]^u[6]^u[3]^u[1]^u[0];
	y[5] = x[299]^x[300]^x[302]^x[304]^x[307]^x[311]^x[312]^x[313]^x[314]^x[315]^x[317]^x[321]^x[323]^x[324]^x[327]^x[329]^u[30]^u[29]^u[27]^u[25]^u[22]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[8]^u[6]^u[5]^u[2]^u[0];
	y[6] = x[300]^x[301]^x[303]^x[305]^x[308]^x[312]^x[313]^x[314]^x[315]^x[316]^x[318]^x[322]^x[324]^x[325]^x[328]^u[29]^u[28]^u[26]^u[24]^u[21]^u[17]^u[16]^u[15]^u[14]^u[13]^u[11]^u[7]^u[5]^u[4]^u[1];
	y[7] = x[301]^x[302]^x[304]^x[306]^x[309]^x[313]^x[314]^x[315]^x[316]^x[317]^x[319]^x[323]^x[325]^x[326]^x[329]^u[28]^u[27]^u[25]^u[23]^u[20]^u[16]^u[15]^u[14]^u[13]^u[12]^u[10]^u[6]^u[4]^u[3]^u[0];
	y[8] = x[302]^x[303]^x[305]^x[307]^x[310]^x[314]^x[315]^x[316]^x[317]^x[318]^x[320]^x[324]^x[326]^x[327]^u[27]^u[26]^u[24]^u[22]^u[19]^u[15]^u[14]^u[13]^u[12]^u[11]^u[9]^u[5]^u[3]^u[2];
	y[9] = x[298]^x[299]^x[300]^x[301]^x[302]^x[303]^x[307]^x[308]^x[310]^x[311]^x[315]^x[317]^x[320]^x[321]^x[323]^x[324]^x[326]^x[328]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[22]^u[21]^u[19]^u[18]^u[14]^u[12]^u[9]^u[8]^u[6]^u[5]^u[3]^u[1];
	y[10] = x[299]^x[300]^x[301]^x[302]^x[303]^x[304]^x[308]^x[309]^x[311]^x[312]^x[316]^x[318]^x[321]^x[322]^x[324]^x[325]^x[327]^x[329]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[21]^u[20]^u[18]^u[17]^u[13]^u[11]^u[8]^u[7]^u[5]^u[4]^u[2]^u[0];
	y[11] = x[300]^x[301]^x[302]^x[303]^x[304]^x[305]^x[309]^x[310]^x[312]^x[313]^x[317]^x[319]^x[322]^x[323]^x[325]^x[326]^x[328]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[20]^u[19]^u[17]^u[16]^u[12]^u[10]^u[7]^u[6]^u[4]^u[3]^u[1];
	y[12] = x[298]^x[299]^x[300]^x[303]^x[305]^x[307]^x[311]^x[313]^x[314]^x[316]^x[319]^x[325]^x[329]^u[31]^u[30]^u[29]^u[26]^u[24]^u[22]^u[18]^u[16]^u[15]^u[13]^u[10]^u[4]^u[0];
	y[13] = x[298]^x[302]^x[307]^x[308]^x[310]^x[312]^x[314]^x[315]^x[316]^x[317]^x[318]^x[319]^x[323]^x[324]^x[325]^x[327]^u[31]^u[27]^u[22]^u[21]^u[19]^u[17]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[6]^u[5]^u[4]^u[2];
	y[14] = x[299]^x[303]^x[308]^x[309]^x[311]^x[313]^x[315]^x[316]^x[317]^x[318]^x[319]^x[320]^x[324]^x[325]^x[326]^x[328]^u[30]^u[26]^u[21]^u[20]^u[18]^u[16]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[5]^u[4]^u[3]^u[1];
	y[15] = x[298]^x[299]^x[301]^x[302]^x[306]^x[307]^x[309]^x[312]^x[314]^x[317]^x[321]^x[323]^x[324]^x[329]^u[31]^u[30]^u[28]^u[27]^u[23]^u[22]^u[20]^u[17]^u[15]^u[12]^u[8]^u[6]^u[5]^u[0];
	y[16] = x[298]^x[301]^x[303]^x[304]^x[306]^x[308]^x[313]^x[315]^x[316]^x[319]^x[320]^x[322]^x[323]^x[326]^x[327]^u[31]^u[28]^u[26]^u[25]^u[23]^u[21]^u[16]^u[14]^u[13]^u[10]^u[9]^u[7]^u[6]^u[3]^u[2];
	y[17] = x[299]^x[302]^x[304]^x[305]^x[307]^x[309]^x[314]^x[316]^x[317]^x[320]^x[321]^x[323]^x[324]^x[327]^x[328]^u[30]^u[27]^u[25]^u[24]^u[22]^u[20]^u[15]^u[13]^u[12]^u[9]^u[8]^u[6]^u[5]^u[2]^u[1];
	y[18] = x[300]^x[303]^x[305]^x[306]^x[308]^x[310]^x[315]^x[317]^x[318]^x[321]^x[322]^x[324]^x[325]^x[328]^x[329]^u[29]^u[26]^u[24]^u[23]^u[21]^u[19]^u[14]^u[12]^u[11]^u[8]^u[7]^u[5]^u[4]^u[1]^u[0];
	y[19] = x[298]^x[299]^x[300]^x[302]^x[309]^x[310]^x[311]^x[320]^x[322]^x[324]^x[327]^x[329]^u[31]^u[30]^u[29]^u[27]^u[20]^u[19]^u[18]^u[9]^u[7]^u[5]^u[2]^u[0];
	y[20] = x[299]^x[300]^x[301]^x[303]^x[310]^x[311]^x[312]^x[321]^x[323]^x[325]^x[328]^u[30]^u[29]^u[28]^u[26]^u[19]^u[18]^u[17]^u[8]^u[6]^u[4]^u[1];
	y[21] = x[300]^x[301]^x[302]^x[304]^x[311]^x[312]^x[313]^x[322]^x[324]^x[326]^x[329]^u[29]^u[28]^u[27]^u[25]^u[18]^u[17]^u[16]^u[7]^u[5]^u[3]^u[0];
	y[22] = x[301]^x[302]^x[303]^x[305]^x[312]^x[313]^x[314]^x[323]^x[325]^x[327]^u[28]^u[27]^u[26]^u[24]^u[17]^u[16]^u[15]^u[6]^u[4]^u[2];
	y[23] = x[302]^x[303]^x[304]^x[306]^x[313]^x[314]^x[315]^x[324]^x[326]^x[328]^u[27]^u[26]^u[25]^u[23]^u[16]^u[15]^u[14]^u[5]^u[3]^u[1];
	y[24] = x[303]^x[304]^x[305]^x[307]^x[314]^x[315]^x[316]^x[325]^x[327]^x[329]^u[26]^u[25]^u[24]^u[22]^u[15]^u[14]^u[13]^u[4]^u[2]^u[0];
	y[25] = x[298]^x[299]^x[300]^x[301]^x[302]^x[305]^x[307]^x[308]^x[310]^x[315]^x[317]^x[318]^x[319]^x[320]^x[323]^x[324]^x[325]^x[327]^x[328]^u[31]^u[30]^u[29]^u[28]^u[27]^u[24]^u[22]^u[21]^u[19]^u[14]^u[12]^u[11]^u[10]^u[9]^u[6]^u[5]^u[4]^u[2]^u[1];
	y[26] = x[299]^x[300]^x[301]^x[302]^x[303]^x[306]^x[308]^x[309]^x[311]^x[316]^x[318]^x[319]^x[320]^x[321]^x[324]^x[325]^x[326]^x[328]^x[329]^u[30]^u[29]^u[28]^u[27]^u[26]^u[23]^u[21]^u[20]^u[18]^u[13]^u[11]^u[10]^u[9]^u[8]^u[5]^u[4]^u[3]^u[1]^u[0];
	y[27] = x[298]^x[299]^x[303]^x[306]^x[309]^x[312]^x[316]^x[317]^x[318]^x[321]^x[322]^x[323]^x[324]^x[329]^u[31]^u[30]^u[26]^u[23]^u[20]^u[17]^u[13]^u[12]^u[11]^u[8]^u[7]^u[6]^u[5]^u[0];
	y[28] = x[298]^x[301]^x[302]^x[306]^x[313]^x[316]^x[317]^x[320]^x[322]^x[326]^x[327]^u[31]^u[28]^u[27]^u[23]^u[16]^u[13]^u[12]^u[9]^u[7]^u[3]^u[2];
	y[29] = x[298]^x[300]^x[301]^x[303]^x[304]^x[306]^x[310]^x[314]^x[316]^x[317]^x[319]^x[320]^x[321]^x[324]^x[325]^x[326]^x[328]^u[31]^u[29]^u[28]^u[26]^u[25]^u[23]^u[19]^u[15]^u[13]^u[12]^u[10]^u[9]^u[8]^u[5]^u[4]^u[3]^u[1];
	y[30] = x[299]^x[301]^x[302]^x[304]^x[305]^x[307]^x[311]^x[315]^x[317]^x[318]^x[320]^x[321]^x[322]^x[325]^x[326]^x[327]^x[329]^u[30]^u[28]^u[27]^u[25]^u[24]^u[22]^u[18]^u[14]^u[12]^u[11]^u[9]^u[8]^u[7]^u[4]^u[3]^u[2]^u[0];
	y[31] = x[298]^x[299]^x[301]^x[303]^x[304]^x[305]^x[307]^x[308]^x[310]^x[312]^x[320]^x[321]^x[322]^x[324]^x[325]^x[328]^u[31]^u[30]^u[28]^u[26]^u[25]^u[24]^u[22]^u[21]^u[19]^u[17]^u[9]^u[8]^u[7]^u[5]^u[4]^u[1];
	y[32] = x[0]^x[298]^x[301]^x[305]^x[307]^x[308]^x[309]^x[310]^x[311]^x[313]^x[316]^x[318]^x[319]^x[320]^x[321]^x[322]^x[324]^x[327]^x[329]^u[31]^u[28]^u[24]^u[22]^u[21]^u[20]^u[19]^u[18]^u[16]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[5]^u[2]^u[0];
	y[33] = x[1]^x[298]^x[300]^x[301]^x[304]^x[307]^x[308]^x[309]^x[311]^x[312]^x[314]^x[316]^x[317]^x[318]^x[321]^x[322]^x[324]^x[326]^x[327]^x[328]^u[31]^u[29]^u[28]^u[25]^u[22]^u[21]^u[20]^u[18]^u[17]^u[15]^u[13]^u[12]^u[11]^u[8]^u[7]^u[5]^u[3]^u[2]^u[1];
	y[34] = x[2]^x[298]^x[300]^x[304]^x[305]^x[306]^x[307]^x[308]^x[309]^x[312]^x[313]^x[315]^x[316]^x[317]^x[320]^x[322]^x[324]^x[326]^x[328]^x[329]^u[31]^u[29]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[17]^u[16]^u[14]^u[13]^u[12]^u[9]^u[7]^u[5]^u[3]^u[1]^u[0];
	y[35] = x[3]^x[299]^x[301]^x[305]^x[306]^x[307]^x[308]^x[309]^x[310]^x[313]^x[314]^x[316]^x[317]^x[318]^x[321]^x[323]^x[325]^x[327]^x[329]^u[30]^u[28]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[16]^u[15]^u[13]^u[12]^u[11]^u[8]^u[6]^u[4]^u[2]^u[0];
	y[36] = x[4]^x[298]^x[299]^x[301]^x[304]^x[308]^x[309]^x[311]^x[314]^x[315]^x[316]^x[317]^x[320]^x[322]^x[323]^x[325]^x[327]^x[328]^u[31]^u[30]^u[28]^u[25]^u[21]^u[20]^u[18]^u[15]^u[14]^u[13]^u[12]^u[9]^u[7]^u[6]^u[4]^u[2]^u[1];
	y[37] = x[5]^x[299]^x[300]^x[302]^x[305]^x[309]^x[310]^x[312]^x[315]^x[316]^x[317]^x[318]^x[321]^x[323]^x[324]^x[326]^x[328]^x[329]^u[30]^u[29]^u[27]^u[24]^u[20]^u[19]^u[17]^u[14]^u[13]^u[12]^u[11]^u[8]^u[6]^u[5]^u[3]^u[1]^u[0];
	y[38] = x[6]^x[298]^x[299]^x[302]^x[303]^x[304]^x[307]^x[311]^x[313]^x[317]^x[320]^x[322]^x[323]^x[326]^x[329]^u[31]^u[30]^u[27]^u[26]^u[25]^u[22]^u[18]^u[16]^u[12]^u[9]^u[7]^u[6]^u[3]^u[0];
	y[39] = x[7]^x[299]^x[300]^x[303]^x[304]^x[305]^x[308]^x[312]^x[314]^x[318]^x[321]^x[323]^x[324]^x[327]^u[30]^u[29]^u[26]^u[25]^u[24]^u[21]^u[17]^u[15]^u[11]^u[8]^u[6]^u[5]^u[2];
	y[40] = x[8]^x[300]^x[301]^x[304]^x[305]^x[306]^x[309]^x[313]^x[315]^x[319]^x[322]^x[324]^x[325]^x[328]^u[29]^u[28]^u[25]^u[24]^u[23]^u[20]^u[16]^u[14]^u[10]^u[7]^u[5]^u[4]^u[1];
	y[41] = x[9]^x[298]^x[299]^x[300]^x[304]^x[305]^x[314]^x[318]^x[319]^x[324]^x[327]^x[329]^u[31]^u[30]^u[29]^u[25]^u[24]^u[15]^u[11]^u[10]^u[5]^u[2]^u[0];
	y[42] = x[10]^x[298]^x[302]^x[304]^x[305]^x[307]^x[310]^x[315]^x[316]^x[318]^x[323]^x[324]^x[326]^x[327]^x[328]^u[31]^u[27]^u[25]^u[24]^u[22]^u[19]^u[14]^u[13]^u[11]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[43] = x[11]^x[299]^x[303]^x[305]^x[306]^x[308]^x[311]^x[316]^x[317]^x[319]^x[324]^x[325]^x[327]^x[328]^x[329]^u[30]^u[26]^u[24]^u[23]^u[21]^u[18]^u[13]^u[12]^u[10]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[44] = x[12]^x[300]^x[304]^x[306]^x[307]^x[309]^x[312]^x[317]^x[318]^x[320]^x[325]^x[326]^x[328]^x[329]^u[29]^u[25]^u[23]^u[22]^u[20]^u[17]^u[12]^u[11]^u[9]^u[4]^u[3]^u[1]^u[0];
	y[45] = x[13]^x[298]^x[299]^x[300]^x[302]^x[304]^x[305]^x[306]^x[308]^x[313]^x[316]^x[320]^x[321]^x[323]^x[324]^x[325]^x[329]^u[31]^u[30]^u[29]^u[27]^u[25]^u[24]^u[23]^u[21]^u[16]^u[13]^u[9]^u[8]^u[6]^u[5]^u[4]^u[0];
	y[46] = x[14]^x[298]^x[302]^x[303]^x[304]^x[305]^x[309]^x[310]^x[314]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[327]^u[31]^u[27]^u[26]^u[25]^u[24]^u[20]^u[19]^u[15]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[2];
	y[47] = x[15]^x[299]^x[303]^x[304]^x[305]^x[306]^x[310]^x[311]^x[315]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[328]^u[30]^u[26]^u[25]^u[24]^u[23]^u[19]^u[18]^u[14]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[1];
	y[48] = x[16]^x[300]^x[304]^x[305]^x[306]^x[307]^x[311]^x[312]^x[316]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[325]^x[329]^u[29]^u[25]^u[24]^u[23]^u[22]^u[18]^u[17]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[0];
	y[49] = x[17]^x[298]^x[299]^x[300]^x[302]^x[304]^x[305]^x[308]^x[310]^x[312]^x[313]^x[316]^x[317]^x[318]^x[321]^x[322]^x[327]^u[31]^u[30]^u[29]^u[27]^u[25]^u[24]^u[21]^u[19]^u[17]^u[16]^u[13]^u[12]^u[11]^u[8]^u[7]^u[2];
	y[50] = x[18]^x[298]^x[302]^x[303]^x[304]^x[305]^x[307]^x[309]^x[310]^x[311]^x[313]^x[314]^x[316]^x[317]^x[320]^x[322]^x[324]^x[325]^x[326]^x[327]^x[328]^u[31]^u[27]^u[26]^u[25]^u[24]^u[22]^u[20]^u[19]^u[18]^u[16]^u[15]^u[13]^u[12]^u[9]^u[7]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[51] = x[19]^x[299]^x[303]^x[304]^x[305]^x[306]^x[308]^x[310]^x[311]^x[312]^x[314]^x[315]^x[317]^x[318]^x[321]^x[323]^x[325]^x[326]^x[327]^x[328]^x[329]^u[30]^u[26]^u[25]^u[24]^u[23]^u[21]^u[19]^u[18]^u[17]^u[15]^u[14]^u[12]^u[11]^u[8]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[52] = x[20]^x[298]^x[299]^x[301]^x[302]^x[305]^x[309]^x[310]^x[311]^x[312]^x[313]^x[315]^x[320]^x[322]^x[323]^x[325]^x[328]^x[329]^u[31]^u[30]^u[28]^u[27]^u[24]^u[20]^u[19]^u[18]^u[17]^u[16]^u[14]^u[9]^u[7]^u[6]^u[4]^u[1]^u[0];
	y[53] = x[21]^x[299]^x[300]^x[302]^x[303]^x[306]^x[310]^x[311]^x[312]^x[313]^x[314]^x[316]^x[321]^x[323]^x[324]^x[326]^x[329]^u[30]^u[29]^u[27]^u[26]^u[23]^u[19]^u[18]^u[17]^u[16]^u[15]^u[13]^u[8]^u[6]^u[5]^u[3]^u[0];
	y[54] = x[22]^x[300]^x[301]^x[303]^x[304]^x[307]^x[311]^x[312]^x[313]^x[314]^x[315]^x[317]^x[322]^x[324]^x[325]^x[327]^u[29]^u[28]^u[26]^u[25]^u[22]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[7]^u[5]^u[4]^u[2];
	y[55] = x[23]^x[298]^x[299]^x[300]^x[305]^x[306]^x[307]^x[308]^x[310]^x[312]^x[313]^x[314]^x[315]^x[319]^x[320]^x[324]^x[327]^x[328]^u[31]^u[30]^u[29]^u[24]^u[23]^u[22]^u[21]^u[19]^u[17]^u[16]^u[15]^u[14]^u[10]^u[9]^u[5]^u[2]^u[1];
	y[56] = x[24]^x[298]^x[302]^x[304]^x[308]^x[309]^x[310]^x[311]^x[313]^x[314]^x[315]^x[318]^x[319]^x[321]^x[323]^x[324]^x[326]^x[327]^x[328]^x[329]^u[31]^u[27]^u[25]^u[21]^u[20]^u[19]^u[18]^u[16]^u[15]^u[14]^u[11]^u[10]^u[8]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[57] = x[25]^x[298]^x[300]^x[301]^x[302]^x[303]^x[304]^x[305]^x[306]^x[307]^x[309]^x[311]^x[312]^x[314]^x[315]^x[318]^x[322]^x[323]^x[326]^x[328]^x[329]^u[31]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[20]^u[18]^u[17]^u[15]^u[14]^u[11]^u[7]^u[6]^u[3]^u[1]^u[0];
	y[58] = x[26]^x[298]^x[300]^x[303]^x[305]^x[308]^x[312]^x[313]^x[315]^x[318]^x[320]^x[325]^x[326]^x[329]^u[31]^u[29]^u[26]^u[24]^u[21]^u[17]^u[16]^u[14]^u[11]^u[9]^u[4]^u[3]^u[0];
	y[59] = x[27]^x[299]^x[301]^x[304]^x[306]^x[309]^x[313]^x[314]^x[316]^x[319]^x[321]^x[326]^x[327]^u[30]^u[28]^u[25]^u[23]^u[20]^u[16]^u[15]^u[13]^u[10]^u[8]^u[3]^u[2];
	y[60] = x[28]^x[298]^x[299]^x[301]^x[304]^x[305]^x[306]^x[314]^x[315]^x[316]^x[317]^x[318]^x[319]^x[322]^x[323]^x[324]^x[325]^x[326]^x[328]^u[31]^u[30]^u[28]^u[25]^u[24]^u[23]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[7]^u[6]^u[5]^u[4]^u[3]^u[1];
	y[61] = x[29]^x[299]^x[300]^x[302]^x[305]^x[306]^x[307]^x[315]^x[316]^x[317]^x[318]^x[319]^x[320]^x[323]^x[324]^x[325]^x[326]^x[327]^x[329]^u[30]^u[29]^u[27]^u[24]^u[23]^u[22]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[6]^u[5]^u[4]^u[3]^u[2]^u[0];
	y[62] = x[30]^x[300]^x[301]^x[303]^x[306]^x[307]^x[308]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[324]^x[325]^x[326]^x[327]^x[328]^u[29]^u[28]^u[26]^u[23]^u[22]^u[21]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[63] = x[31]^x[301]^x[302]^x[304]^x[307]^x[308]^x[309]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[325]^x[326]^x[327]^x[328]^x[329]^u[28]^u[27]^u[25]^u[22]^u[21]^u[20]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[64] = x[32]^x[298]^x[299]^x[300]^x[301]^x[303]^x[304]^x[305]^x[306]^x[307]^x[308]^x[309]^x[316]^x[321]^x[322]^x[324]^x[325]^x[328]^x[329]^u[31]^u[30]^u[29]^u[28]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[13]^u[8]^u[7]^u[5]^u[4]^u[1]^u[0];
	y[65] = x[33]^x[298]^x[305]^x[308]^x[309]^x[316]^x[317]^x[318]^x[319]^x[320]^x[322]^x[324]^x[327]^x[329]^u[31]^u[24]^u[21]^u[20]^u[13]^u[12]^u[11]^u[10]^u[9]^u[7]^u[5]^u[2]^u[0];
	y[66] = x[34]^x[299]^x[306]^x[309]^x[310]^x[317]^x[318]^x[319]^x[320]^x[321]^x[323]^x[325]^x[328]^u[30]^u[23]^u[20]^u[19]^u[12]^u[11]^u[10]^u[9]^u[8]^u[6]^u[4]^u[1];
	y[67] = x[35]^x[298]^x[299]^x[301]^x[302]^x[304]^x[306]^x[311]^x[316]^x[321]^x[322]^x[323]^x[325]^x[327]^x[329]^u[31]^u[30]^u[28]^u[27]^u[25]^u[23]^u[18]^u[13]^u[8]^u[7]^u[6]^u[4]^u[2]^u[0];
	y[68] = x[36]^x[299]^x[300]^x[302]^x[303]^x[305]^x[307]^x[312]^x[317]^x[322]^x[323]^x[324]^x[326]^x[328]^u[30]^u[29]^u[27]^u[26]^u[24]^u[22]^u[17]^u[12]^u[7]^u[6]^u[5]^u[3]^u[1];
	y[69] = x[37]^x[298]^x[299]^x[302]^x[303]^x[307]^x[308]^x[310]^x[313]^x[316]^x[319]^x[320]^x[326]^x[329]^u[31]^u[30]^u[27]^u[26]^u[22]^u[21]^u[19]^u[16]^u[13]^u[10]^u[9]^u[3]^u[0];
	y[70] = x[38]^x[299]^x[300]^x[303]^x[304]^x[308]^x[309]^x[311]^x[314]^x[317]^x[320]^x[321]^x[327]^u[30]^u[29]^u[26]^u[25]^u[21]^u[20]^u[18]^u[15]^u[12]^u[9]^u[8]^u[2];
	y[71] = x[39]^x[298]^x[299]^x[302]^x[305]^x[306]^x[307]^x[309]^x[312]^x[315]^x[316]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[325]^x[326]^x[327]^x[328]^u[31]^u[30]^u[27]^u[24]^u[23]^u[22]^u[20]^u[17]^u[14]^u[13]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[72] = x[40]^x[298]^x[301]^x[302]^x[303]^x[304]^x[308]^x[313]^x[317]^x[318]^x[319]^x[321]^x[322]^x[328]^x[329]^u[31]^u[28]^u[27]^u[26]^u[25]^u[21]^u[16]^u[12]^u[11]^u[10]^u[8]^u[7]^u[1]^u[0];
	y[73] = x[41]^x[299]^x[302]^x[303]^x[304]^x[305]^x[309]^x[314]^x[318]^x[319]^x[320]^x[322]^x[323]^x[329]^u[30]^u[27]^u[26]^u[25]^u[24]^u[20]^u[15]^u[11]^u[10]^u[9]^u[7]^u[6]^u[0];
	y[74] = x[42]^x[298]^x[299]^x[301]^x[302]^x[303]^x[305]^x[307]^x[315]^x[316]^x[318]^x[321]^x[325]^x[326]^x[327]^u[31]^u[30]^u[28]^u[27]^u[26]^u[24]^u[22]^u[14]^u[13]^u[11]^u[8]^u[4]^u[3]^u[2];
	y[75] = x[43]^x[299]^x[300]^x[302]^x[303]^x[304]^x[306]^x[308]^x[316]^x[317]^x[319]^x[322]^x[326]^x[327]^x[328]^u[30]^u[29]^u[27]^u[26]^u[25]^u[23]^u[21]^u[13]^u[12]^u[10]^u[7]^u[3]^u[2]^u[1];
	y[76] = x[44]^x[300]^x[301]^x[303]^x[304]^x[305]^x[307]^x[309]^x[317]^x[318]^x[320]^x[323]^x[327]^x[328]^x[329]^u[29]^u[28]^u[26]^u[25]^u[24]^u[22]^u[20]^u[12]^u[11]^u[9]^u[6]^u[2]^u[1]^u[0];
	y[77] = x[45]^x[298]^x[299]^x[300]^x[305]^x[307]^x[308]^x[316]^x[320]^x[321]^x[323]^x[325]^x[326]^x[327]^x[328]^x[329]^u[31]^u[30]^u[29]^u[24]^u[22]^u[21]^u[13]^u[9]^u[8]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[78] = x[46]^x[299]^x[300]^x[301]^x[306]^x[308]^x[309]^x[317]^x[321]^x[322]^x[324]^x[326]^x[327]^x[328]^x[329]^u[30]^u[29]^u[28]^u[23]^u[21]^u[20]^u[12]^u[8]^u[7]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[79] = x[47]^x[298]^x[299]^x[304]^x[306]^x[309]^x[316]^x[319]^x[320]^x[322]^x[324]^x[326]^x[328]^x[329]^u[31]^u[30]^u[25]^u[23]^u[20]^u[13]^u[10]^u[9]^u[7]^u[5]^u[3]^u[1]^u[0];
	y[80] = x[48]^x[298]^x[301]^x[302]^x[304]^x[305]^x[306]^x[316]^x[317]^x[318]^x[319]^x[321]^x[324]^x[326]^x[329]^u[31]^u[28]^u[27]^u[25]^u[24]^u[23]^u[13]^u[12]^u[11]^u[10]^u[8]^u[5]^u[3]^u[0];
	y[81] = x[49]^x[299]^x[302]^x[303]^x[305]^x[306]^x[307]^x[317]^x[318]^x[319]^x[320]^x[322]^x[325]^x[327]^u[30]^u[27]^u[26]^u[24]^u[23]^u[22]^u[12]^u[11]^u[10]^u[9]^u[7]^u[4]^u[2];
	y[82] = x[50]^x[298]^x[299]^x[301]^x[302]^x[303]^x[308]^x[310]^x[316]^x[321]^x[324]^x[325]^x[327]^x[328]^u[31]^u[30]^u[28]^u[27]^u[26]^u[21]^u[19]^u[13]^u[8]^u[5]^u[4]^u[2]^u[1];
	y[83] = x[51]^x[298]^x[301]^x[303]^x[306]^x[307]^x[309]^x[310]^x[311]^x[316]^x[317]^x[318]^x[319]^x[320]^x[322]^x[323]^x[324]^x[327]^x[328]^x[329]^u[31]^u[28]^u[26]^u[23]^u[22]^u[20]^u[19]^u[18]^u[13]^u[12]^u[11]^u[10]^u[9]^u[7]^u[6]^u[5]^u[2]^u[1]^u[0];
	y[84] = x[52]^x[299]^x[302]^x[304]^x[307]^x[308]^x[310]^x[311]^x[312]^x[317]^x[318]^x[319]^x[320]^x[321]^x[323]^x[324]^x[325]^x[328]^x[329]^u[30]^u[27]^u[25]^u[22]^u[21]^u[19]^u[18]^u[17]^u[12]^u[11]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4]^u[1]^u[0];
	y[85] = x[53]^x[298]^x[299]^x[301]^x[302]^x[303]^x[304]^x[305]^x[306]^x[307]^x[308]^x[309]^x[310]^x[311]^x[312]^x[313]^x[316]^x[321]^x[322]^x[323]^x[327]^x[329]^u[31]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[13]^u[8]^u[7]^u[6]^u[2]^u[0];
	y[86] = x[54]^x[298]^x[301]^x[303]^x[305]^x[308]^x[309]^x[311]^x[312]^x[313]^x[314]^x[316]^x[317]^x[318]^x[319]^x[320]^x[322]^x[325]^x[326]^x[327]^x[328]^u[31]^u[28]^u[26]^u[24]^u[21]^u[20]^u[18]^u[17]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[9]^u[7]^u[4]^u[3]^u[2]^u[1];
	y[87] = x[55]^x[299]^x[302]^x[304]^x[306]^x[309]^x[310]^x[312]^x[313]^x[314]^x[315]^x[317]^x[318]^x[319]^x[320]^x[321]^x[323]^x[326]^x[327]^x[328]^x[329]^u[30]^u[27]^u[25]^u[23]^u[20]^u[19]^u[17]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[8]^u[6]^u[3]^u[2]^u[1]^u[0];
	y[88] = x[56]^x[300]^x[303]^x[305]^x[307]^x[310]^x[311]^x[313]^x[314]^x[315]^x[316]^x[318]^x[319]^x[320]^x[321]^x[322]^x[324]^x[327]^x[328]^x[329]^u[29]^u[26]^u[24]^u[22]^u[19]^u[18]^u[16]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[5]^u[2]^u[1]^u[0];
	y[89] = x[57]^x[298]^x[299]^x[300]^x[302]^x[307]^x[308]^x[310]^x[311]^x[312]^x[314]^x[315]^x[317]^x[318]^x[321]^x[322]^x[324]^x[326]^x[327]^x[328]^x[329]^u[31]^u[30]^u[29]^u[27]^u[22]^u[21]^u[19]^u[18]^u[17]^u[15]^u[14]^u[12]^u[11]^u[8]^u[7]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[90] = x[58]^x[299]^x[300]^x[301]^x[303]^x[308]^x[309]^x[311]^x[312]^x[313]^x[315]^x[316]^x[318]^x[319]^x[322]^x[323]^x[325]^x[327]^x[328]^x[329]^u[30]^u[29]^u[28]^u[26]^u[21]^u[20]^u[18]^u[17]^u[16]^u[14]^u[13]^u[11]^u[10]^u[7]^u[6]^u[4]^u[2]^u[1]^u[0];
	y[91] = x[59]^x[298]^x[299]^x[306]^x[307]^x[309]^x[312]^x[313]^x[314]^x[317]^x[318]^x[325]^x[327]^x[328]^x[329]^u[31]^u[30]^u[23]^u[22]^u[20]^u[17]^u[16]^u[15]^u[12]^u[11]^u[4]^u[2]^u[1]^u[0];
	y[92] = x[60]^x[298]^x[301]^x[302]^x[304]^x[306]^x[308]^x[313]^x[314]^x[315]^x[316]^x[320]^x[323]^x[324]^x[325]^x[327]^x[328]^x[329]^u[31]^u[28]^u[27]^u[25]^u[23]^u[21]^u[16]^u[15]^u[14]^u[13]^u[9]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[93] = x[61]^x[298]^x[300]^x[301]^x[303]^x[304]^x[305]^x[306]^x[309]^x[310]^x[314]^x[315]^x[317]^x[318]^x[319]^x[320]^x[321]^x[323]^x[327]^x[328]^x[329]^u[31]^u[29]^u[28]^u[26]^u[25]^u[24]^u[23]^u[20]^u[19]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[8]^u[6]^u[2]^u[1]^u[0];
	y[94] = x[62]^x[299]^x[301]^x[302]^x[304]^x[305]^x[306]^x[307]^x[310]^x[311]^x[315]^x[316]^x[318]^x[319]^x[320]^x[321]^x[322]^x[324]^x[328]^x[329]^u[30]^u[28]^u[27]^u[25]^u[24]^u[23]^u[22]^u[19]^u[18]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[5]^u[1]^u[0];
	y[95] = x[63]^x[298]^x[299]^x[301]^x[303]^x[304]^x[305]^x[308]^x[310]^x[311]^x[312]^x[317]^x[318]^x[321]^x[322]^x[324]^x[326]^x[327]^x[329]^u[31]^u[30]^u[28]^u[26]^u[25]^u[24]^u[21]^u[19]^u[18]^u[17]^u[12]^u[11]^u[8]^u[7]^u[5]^u[3]^u[2]^u[0];
	y[96] = x[64]^x[298]^x[301]^x[305]^x[307]^x[309]^x[310]^x[311]^x[312]^x[313]^x[316]^x[320]^x[322]^x[324]^x[326]^x[328]^u[31]^u[28]^u[24]^u[22]^u[20]^u[19]^u[18]^u[17]^u[16]^u[13]^u[9]^u[7]^u[5]^u[3]^u[1];
	y[97] = x[65]^x[298]^x[300]^x[301]^x[304]^x[307]^x[308]^x[311]^x[312]^x[313]^x[314]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[324]^x[326]^x[329]^u[31]^u[29]^u[28]^u[25]^u[22]^u[21]^u[18]^u[17]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[5]^u[3]^u[0];
	y[98] = x[66]^x[298]^x[300]^x[304]^x[305]^x[306]^x[307]^x[308]^x[309]^x[310]^x[312]^x[313]^x[314]^x[315]^x[316]^x[317]^x[321]^x[322]^x[323]^x[324]^x[326]^u[31]^u[29]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[17]^u[16]^u[15]^u[14]^u[13]^u[12]^u[8]^u[7]^u[6]^u[5]^u[3];
	y[99] = x[67]^x[299]^x[301]^x[305]^x[306]^x[307]^x[308]^x[309]^x[310]^x[311]^x[313]^x[314]^x[315]^x[316]^x[317]^x[318]^x[322]^x[323]^x[324]^x[325]^x[327]^u[30]^u[28]^u[24]^u[23]^u[22]^u[21]^u[20]^u[19]^u[18]^u[16]^u[15]^u[14]^u[13]^u[12]^u[11]^u[7]^u[6]^u[5]^u[4]^u[2];
	y[100] = x[68]^x[298]^x[299]^x[301]^x[304]^x[308]^x[309]^x[311]^x[312]^x[314]^x[315]^x[317]^x[320]^x[327]^x[328]^u[31]^u[30]^u[28]^u[25]^u[21]^u[20]^u[18]^u[17]^u[15]^u[14]^u[12]^u[9]^u[2]^u[1];
	y[101] = x[69]^x[299]^x[300]^x[302]^x[305]^x[309]^x[310]^x[312]^x[313]^x[315]^x[316]^x[318]^x[321]^x[328]^x[329]^u[30]^u[29]^u[27]^u[24]^u[20]^u[19]^u[17]^u[16]^u[14]^u[13]^u[11]^u[8]^u[1]^u[0];
	y[102] = x[70]^x[300]^x[301]^x[303]^x[306]^x[310]^x[311]^x[313]^x[314]^x[316]^x[317]^x[319]^x[322]^x[329]^u[29]^u[28]^u[26]^u[23]^u[19]^u[18]^u[16]^u[15]^u[13]^u[12]^u[10]^u[7]^u[0];
	y[103] = x[71]^x[301]^x[302]^x[304]^x[307]^x[311]^x[312]^x[314]^x[315]^x[317]^x[318]^x[320]^x[323]^u[28]^u[27]^u[25]^u[22]^u[18]^u[17]^u[15]^u[14]^u[12]^u[11]^u[9]^u[6];
	y[104] = x[72]^x[302]^x[303]^x[305]^x[308]^x[312]^x[313]^x[315]^x[316]^x[318]^x[319]^x[321]^x[324]^u[27]^u[26]^u[24]^u[21]^u[17]^u[16]^u[14]^u[13]^u[11]^u[10]^u[8]^u[5];
	y[105] = x[73]^x[303]^x[304]^x[306]^x[309]^x[313]^x[314]^x[316]^x[317]^x[319]^x[320]^x[322]^x[325]^u[26]^u[25]^u[23]^u[20]^u[16]^u[15]^u[13]^u[12]^u[10]^u[9]^u[7]^u[4];
	y[106] = x[74]^x[298]^x[299]^x[300]^x[301]^x[302]^x[305]^x[306]^x[314]^x[315]^x[316]^x[317]^x[319]^x[321]^x[324]^x[325]^x[327]^u[31]^u[30]^u[29]^u[28]^u[27]^u[24]^u[23]^u[15]^u[14]^u[13]^u[12]^u[10]^u[8]^u[5]^u[4]^u[2];
	y[107] = x[75]^x[298]^x[303]^x[304]^x[310]^x[315]^x[317]^x[319]^x[322]^x[323]^x[324]^x[327]^x[328]^u[31]^u[26]^u[25]^u[19]^u[14]^u[12]^u[10]^u[7]^u[6]^u[5]^u[2]^u[1];
	y[108] = x[76]^x[299]^x[304]^x[305]^x[311]^x[316]^x[318]^x[320]^x[323]^x[324]^x[325]^x[328]^x[329]^u[30]^u[25]^u[24]^u[18]^u[13]^u[11]^u[9]^u[6]^u[5]^u[4]^u[1]^u[0];
	y[109] = x[77]^x[298]^x[299]^x[301]^x[302]^x[304]^x[305]^x[307]^x[310]^x[312]^x[316]^x[317]^x[318]^x[320]^x[321]^x[323]^x[327]^x[329]^u[31]^u[30]^u[28]^u[27]^u[25]^u[24]^u[22]^u[19]^u[17]^u[13]^u[12]^u[11]^u[9]^u[8]^u[6]^u[2]^u[0];
	y[110] = x[78]^x[299]^x[300]^x[302]^x[303]^x[305]^x[306]^x[308]^x[311]^x[313]^x[317]^x[318]^x[319]^x[321]^x[322]^x[324]^x[328]^u[30]^u[29]^u[27]^u[26]^u[24]^u[23]^u[21]^u[18]^u[16]^u[12]^u[11]^u[10]^u[8]^u[7]^u[5]^u[1];
	y[111] = x[79]^x[298]^x[299]^x[302]^x[303]^x[309]^x[310]^x[312]^x[314]^x[316]^x[322]^x[324]^x[326]^x[327]^x[329]^u[31]^u[30]^u[27]^u[26]^u[20]^u[19]^u[17]^u[15]^u[13]^u[7]^u[5]^u[3]^u[2]^u[0];
	y[112] = x[80]^x[299]^x[300]^x[303]^x[304]^x[310]^x[311]^x[313]^x[315]^x[317]^x[323]^x[325]^x[327]^x[328]^u[30]^u[29]^u[26]^u[25]^u[19]^u[18]^u[16]^u[14]^u[12]^u[6]^u[4]^u[2]^u[1];
	y[113] = x[81]^x[300]^x[301]^x[304]^x[305]^x[311]^x[312]^x[314]^x[316]^x[318]^x[324]^x[326]^x[328]^x[329]^u[29]^u[28]^u[25]^u[24]^u[18]^u[17]^u[15]^u[13]^u[11]^u[5]^u[3]^u[1]^u[0];
	y[114] = x[82]^x[298]^x[299]^x[300]^x[304]^x[305]^x[307]^x[310]^x[312]^x[313]^x[315]^x[316]^x[317]^x[318]^x[320]^x[323]^x[324]^x[326]^x[329]^u[31]^u[30]^u[29]^u[25]^u[24]^u[22]^u[19]^u[17]^u[16]^u[14]^u[13]^u[12]^u[11]^u[9]^u[6]^u[5]^u[3]^u[0];
	y[115] = x[83]^x[299]^x[300]^x[301]^x[305]^x[306]^x[308]^x[311]^x[313]^x[314]^x[316]^x[317]^x[318]^x[319]^x[321]^x[324]^x[325]^x[327]^u[30]^u[29]^u[28]^u[24]^u[23]^u[21]^u[18]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[8]^u[5]^u[4]^u[2];
	y[116] = x[84]^x[300]^x[301]^x[302]^x[306]^x[307]^x[309]^x[312]^x[314]^x[315]^x[317]^x[318]^x[319]^x[320]^x[322]^x[325]^x[326]^x[328]^u[29]^u[28]^u[27]^u[23]^u[22]^u[20]^u[17]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[7]^u[4]^u[3]^u[1];
	y[117] = x[85]^x[298]^x[299]^x[300]^x[303]^x[304]^x[306]^x[308]^x[313]^x[315]^x[321]^x[324]^x[325]^x[329]^u[31]^u[30]^u[29]^u[26]^u[25]^u[23]^u[21]^u[16]^u[14]^u[8]^u[5]^u[4]^u[0];
	y[118] = x[86]^x[299]^x[300]^x[301]^x[304]^x[305]^x[307]^x[309]^x[314]^x[316]^x[322]^x[325]^x[326]^u[30]^u[29]^u[28]^u[25]^u[24]^u[22]^u[20]^u[15]^u[13]^u[7]^u[4]^u[3];
	y[119] = x[87]^x[300]^x[301]^x[302]^x[305]^x[306]^x[308]^x[310]^x[315]^x[317]^x[323]^x[326]^x[327]^u[29]^u[28]^u[27]^u[24]^u[23]^u[21]^u[19]^u[14]^u[12]^u[6]^u[3]^u[2];
	y[120] = x[88]^x[301]^x[302]^x[303]^x[306]^x[307]^x[309]^x[311]^x[316]^x[318]^x[324]^x[327]^x[328]^u[28]^u[27]^u[26]^u[23]^u[22]^u[20]^u[18]^u[13]^u[11]^u[5]^u[2]^u[1];
	y[121] = x[89]^x[302]^x[303]^x[304]^x[307]^x[308]^x[310]^x[312]^x[317]^x[319]^x[325]^x[328]^x[329]^u[27]^u[26]^u[25]^u[22]^u[21]^u[19]^u[17]^u[12]^u[10]^u[4]^u[1]^u[0];
	y[122] = x[90]^x[303]^x[304]^x[305]^x[308]^x[309]^x[311]^x[313]^x[318]^x[320]^x[326]^x[329]^u[26]^u[25]^u[24]^u[21]^u[20]^u[18]^u[16]^u[11]^u[9]^u[3]^u[0];
	y[123] = x[91]^x[304]^x[305]^x[306]^x[309]^x[310]^x[312]^x[314]^x[319]^x[321]^x[327]^u[25]^u[24]^u[23]^u[20]^u[19]^u[17]^u[15]^u[10]^u[8]^u[2];
	y[124] = x[92]^x[298]^x[299]^x[300]^x[301]^x[302]^x[304]^x[305]^x[311]^x[313]^x[315]^x[316]^x[318]^x[319]^x[322]^x[323]^x[324]^x[325]^x[326]^x[327]^x[328]^u[31]^u[30]^u[29]^u[28]^u[27]^u[25]^u[24]^u[18]^u[16]^u[14]^u[13]^u[11]^u[10]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[125] = x[93]^x[299]^x[300]^x[301]^x[302]^x[303]^x[305]^x[306]^x[312]^x[314]^x[316]^x[317]^x[319]^x[320]^x[323]^x[324]^x[325]^x[326]^x[327]^x[328]^x[329]^u[30]^u[29]^u[28]^u[27]^u[26]^u[24]^u[23]^u[17]^u[15]^u[13]^u[12]^u[10]^u[9]^u[6]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[126] = x[94]^x[300]^x[301]^x[302]^x[303]^x[304]^x[306]^x[307]^x[313]^x[315]^x[317]^x[318]^x[320]^x[321]^x[324]^x[325]^x[326]^x[327]^x[328]^x[329]^u[29]^u[28]^u[27]^u[26]^u[25]^u[23]^u[22]^u[16]^u[14]^u[12]^u[11]^u[9]^u[8]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[127] = x[95]^x[298]^x[299]^x[300]^x[303]^x[305]^x[306]^x[308]^x[310]^x[314]^x[320]^x[321]^x[322]^x[323]^x[324]^x[328]^x[329]^u[31]^u[30]^u[29]^u[26]^u[24]^u[23]^u[21]^u[19]^u[15]^u[9]^u[8]^u[7]^u[6]^u[5]^u[1]^u[0];
	y[128] = x[96]^x[299]^x[300]^x[301]^x[304]^x[306]^x[307]^x[309]^x[311]^x[315]^x[321]^x[322]^x[323]^x[324]^x[325]^x[329]^u[30]^u[29]^u[28]^u[25]^u[23]^u[22]^u[20]^u[18]^u[14]^u[8]^u[7]^u[6]^u[5]^u[4]^u[0];
	y[129] = x[97]^x[300]^x[301]^x[302]^x[305]^x[307]^x[308]^x[310]^x[312]^x[316]^x[322]^x[323]^x[324]^x[325]^x[326]^u[29]^u[28]^u[27]^u[24]^u[22]^u[21]^u[19]^u[17]^u[13]^u[7]^u[6]^u[5]^u[4]^u[3];
	y[130] = x[98]^x[298]^x[299]^x[300]^x[303]^x[304]^x[307]^x[308]^x[309]^x[310]^x[311]^x[313]^x[316]^x[317]^x[318]^x[319]^x[320]^u[31]^u[30]^u[29]^u[26]^u[25]^u[22]^u[21]^u[20]^u[19]^u[18]^u[16]^u[13]^u[12]^u[11]^u[10]^u[9];
	y[131] = x[99]^x[298]^x[302]^x[305]^x[306]^x[307]^x[308]^x[309]^x[311]^x[312]^x[314]^x[316]^x[317]^x[321]^x[323]^x[324]^x[325]^x[326]^x[327]^u[31]^u[27]^u[24]^u[23]^u[22]^u[21]^u[20]^u[18]^u[17]^u[15]^u[13]^u[12]^u[8]^u[6]^u[5]^u[4]^u[3]^u[2];
	y[132] = x[100]^x[299]^x[303]^x[306]^x[307]^x[308]^x[309]^x[310]^x[312]^x[313]^x[315]^x[317]^x[318]^x[322]^x[324]^x[325]^x[326]^x[327]^x[328]^u[30]^u[26]^u[23]^u[22]^u[21]^u[20]^u[19]^u[17]^u[16]^u[14]^u[12]^u[11]^u[7]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[133] = x[101]^x[300]^x[304]^x[307]^x[308]^x[309]^x[310]^x[311]^x[313]^x[314]^x[316]^x[318]^x[319]^x[323]^x[325]^x[326]^x[327]^x[328]^x[329]^u[29]^u[25]^u[22]^u[21]^u[20]^u[19]^u[18]^u[16]^u[15]^u[13]^u[11]^u[10]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[134] = x[102]^x[298]^x[299]^x[300]^x[302]^x[304]^x[305]^x[306]^x[307]^x[308]^x[309]^x[311]^x[312]^x[314]^x[315]^x[316]^x[317]^x[318]^x[323]^x[325]^x[328]^x[329]^u[31]^u[30]^u[29]^u[27]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[18]^u[17]^u[15]^u[14]^u[13]^u[12]^u[11]^u[6]^u[4]^u[1]^u[0];
	y[135] = x[103]^x[298]^x[302]^x[303]^x[304]^x[305]^x[308]^x[309]^x[312]^x[313]^x[315]^x[317]^x[320]^x[323]^x[325]^x[327]^x[329]^u[31]^u[27]^u[26]^u[25]^u[24]^u[21]^u[20]^u[17]^u[16]^u[14]^u[12]^u[9]^u[6]^u[4]^u[2]^u[0];
	y[136] = x[104]^x[299]^x[303]^x[304]^x[305]^x[306]^x[309]^x[310]^x[313]^x[314]^x[316]^x[318]^x[321]^x[324]^x[326]^x[328]^u[30]^u[26]^u[25]^u[24]^u[23]^u[20]^u[19]^u[16]^u[15]^u[13]^u[11]^u[8]^u[5]^u[3]^u[1];
	y[137] = x[105]^x[298]^x[299]^x[301]^x[302]^x[305]^x[311]^x[314]^x[315]^x[316]^x[317]^x[318]^x[320]^x[322]^x[323]^x[324]^x[326]^x[329]^u[31]^u[30]^u[28]^u[27]^u[24]^u[18]^u[15]^u[14]^u[13]^u[12]^u[11]^u[9]^u[7]^u[6]^u[5]^u[3]^u[0];
	y[138] = x[106]^x[299]^x[300]^x[302]^x[303]^x[306]^x[312]^x[315]^x[316]^x[317]^x[318]^x[319]^x[321]^x[323]^x[324]^x[325]^x[327]^u[30]^u[29]^u[27]^u[26]^u[23]^u[17]^u[14]^u[13]^u[12]^u[11]^u[10]^u[8]^u[6]^u[5]^u[4]^u[2];
	y[139] = x[107]^x[298]^x[299]^x[302]^x[303]^x[306]^x[310]^x[313]^x[317]^x[322]^x[323]^x[327]^x[328]^u[31]^u[30]^u[27]^u[26]^u[23]^u[19]^u[16]^u[12]^u[7]^u[6]^u[2]^u[1];
	y[140] = x[108]^x[299]^x[300]^x[303]^x[304]^x[307]^x[311]^x[314]^x[318]^x[323]^x[324]^x[328]^x[329]^u[30]^u[29]^u[26]^u[25]^u[22]^u[18]^u[15]^u[11]^u[6]^u[5]^u[1]^u[0];
	y[141] = x[109]^x[298]^x[299]^x[302]^x[305]^x[306]^x[307]^x[308]^x[310]^x[312]^x[315]^x[316]^x[318]^x[320]^x[323]^x[326]^x[327]^x[329]^u[31]^u[30]^u[27]^u[24]^u[23]^u[22]^u[21]^u[19]^u[17]^u[14]^u[13]^u[11]^u[9]^u[6]^u[3]^u[2]^u[0];
	y[142] = x[110]^x[299]^x[300]^x[303]^x[306]^x[307]^x[308]^x[309]^x[311]^x[313]^x[316]^x[317]^x[319]^x[321]^x[324]^x[327]^x[328]^u[30]^u[29]^u[26]^u[23]^u[22]^u[21]^u[20]^u[18]^u[16]^u[13]^u[12]^u[10]^u[8]^u[5]^u[2]^u[1];
	y[143] = x[111]^x[298]^x[299]^x[302]^x[306]^x[308]^x[309]^x[312]^x[314]^x[316]^x[317]^x[319]^x[322]^x[323]^x[324]^x[326]^x[327]^x[328]^x[329]^u[31]^u[30]^u[27]^u[23]^u[21]^u[20]^u[17]^u[15]^u[13]^u[12]^u[10]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[144] = x[112]^x[299]^x[300]^x[303]^x[307]^x[309]^x[310]^x[313]^x[315]^x[317]^x[318]^x[320]^x[323]^x[324]^x[325]^x[327]^x[328]^x[329]^u[30]^u[29]^u[26]^u[22]^u[20]^u[19]^u[16]^u[14]^u[12]^u[11]^u[9]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[145] = x[113]^x[298]^x[299]^x[302]^x[306]^x[307]^x[308]^x[311]^x[314]^x[320]^x[321]^x[323]^x[327]^x[328]^x[329]^u[31]^u[30]^u[27]^u[23]^u[22]^u[21]^u[18]^u[15]^u[9]^u[8]^u[6]^u[2]^u[1]^u[0];
	y[146] = x[114]^x[298]^x[301]^x[302]^x[303]^x[304]^x[306]^x[308]^x[309]^x[310]^x[312]^x[315]^x[316]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[325]^x[326]^x[327]^x[328]^x[329]^u[31]^u[28]^u[27]^u[26]^u[25]^u[23]^u[21]^u[20]^u[19]^u[17]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[147] = x[115]^x[299]^x[302]^x[303]^x[304]^x[305]^x[307]^x[309]^x[310]^x[311]^x[313]^x[316]^x[317]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[326]^x[327]^x[328]^x[329]^u[30]^u[27]^u[26]^u[25]^u[24]^u[22]^u[20]^u[19]^u[18]^u[16]^u[13]^u[12]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[148] = x[116]^x[298]^x[299]^x[301]^x[302]^x[303]^x[305]^x[307]^x[308]^x[311]^x[312]^x[314]^x[316]^x[317]^x[319]^x[321]^x[322]^x[326]^x[328]^x[329]^u[31]^u[30]^u[28]^u[27]^u[26]^u[24]^u[22]^u[21]^u[18]^u[17]^u[15]^u[13]^u[12]^u[10]^u[8]^u[7]^u[3]^u[1]^u[0];
	y[149] = x[117]^x[299]^x[300]^x[302]^x[303]^x[304]^x[306]^x[308]^x[309]^x[312]^x[313]^x[315]^x[317]^x[318]^x[320]^x[322]^x[323]^x[327]^x[329]^u[30]^u[29]^u[27]^u[26]^u[25]^u[23]^u[21]^u[20]^u[17]^u[16]^u[14]^u[12]^u[11]^u[9]^u[7]^u[6]^u[2]^u[0];
	y[150] = x[118]^x[300]^x[301]^x[303]^x[304]^x[305]^x[307]^x[309]^x[310]^x[313]^x[314]^x[316]^x[318]^x[319]^x[321]^x[323]^x[324]^x[328]^u[29]^u[28]^u[26]^u[25]^u[24]^u[22]^u[20]^u[19]^u[16]^u[15]^u[13]^u[11]^u[10]^u[8]^u[6]^u[5]^u[1];
	y[151] = x[119]^x[301]^x[302]^x[304]^x[305]^x[306]^x[308]^x[310]^x[311]^x[314]^x[315]^x[317]^x[319]^x[320]^x[322]^x[324]^x[325]^x[329]^u[28]^u[27]^u[25]^u[24]^u[23]^u[21]^u[19]^u[18]^u[15]^u[14]^u[12]^u[10]^u[9]^u[7]^u[5]^u[4]^u[0];
	y[152] = x[120]^x[298]^x[299]^x[300]^x[301]^x[303]^x[304]^x[305]^x[309]^x[310]^x[311]^x[312]^x[315]^x[319]^x[321]^x[324]^x[327]^u[31]^u[30]^u[29]^u[28]^u[26]^u[25]^u[24]^u[20]^u[19]^u[18]^u[17]^u[14]^u[10]^u[8]^u[5]^u[2];
	y[153] = x[121]^x[299]^x[300]^x[301]^x[302]^x[304]^x[305]^x[306]^x[310]^x[311]^x[312]^x[313]^x[316]^x[320]^x[322]^x[325]^x[328]^u[30]^u[29]^u[28]^u[27]^u[25]^u[24]^u[23]^u[19]^u[18]^u[17]^u[16]^u[13]^u[9]^u[7]^u[4]^u[1];
	y[154] = x[122]^x[298]^x[299]^x[303]^x[304]^x[305]^x[310]^x[311]^x[312]^x[313]^x[314]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[324]^x[325]^x[327]^x[329]^u[31]^u[30]^u[26]^u[25]^u[24]^u[19]^u[18]^u[17]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[5]^u[4]^u[2]^u[0];
	y[155] = x[123]^x[299]^x[300]^x[304]^x[305]^x[306]^x[311]^x[312]^x[313]^x[314]^x[315]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[325]^x[326]^x[328]^u[30]^u[29]^u[25]^u[24]^u[23]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[4]^u[3]^u[1];
	y[156] = x[124]^x[300]^x[301]^x[305]^x[306]^x[307]^x[312]^x[313]^x[314]^x[315]^x[316]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[326]^x[327]^x[329]^u[29]^u[28]^u[24]^u[23]^u[22]^u[17]^u[16]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[3]^u[2]^u[0];
	y[157] = x[125]^x[298]^x[299]^x[300]^x[304]^x[308]^x[310]^x[313]^x[314]^x[315]^x[317]^x[318]^x[321]^x[322]^x[325]^x[326]^x[328]^u[31]^u[30]^u[29]^u[25]^u[21]^u[19]^u[16]^u[15]^u[14]^u[12]^u[11]^u[8]^u[7]^u[4]^u[3]^u[1];
	y[158] = x[126]^x[299]^x[300]^x[301]^x[305]^x[309]^x[311]^x[314]^x[315]^x[316]^x[318]^x[319]^x[322]^x[323]^x[326]^x[327]^x[329]^u[30]^u[29]^u[28]^u[24]^u[20]^u[18]^u[15]^u[14]^u[13]^u[11]^u[10]^u[7]^u[6]^u[3]^u[2]^u[0];
	y[159] = x[127]^x[298]^x[299]^x[304]^x[307]^x[312]^x[315]^x[317]^x[318]^x[325]^x[326]^x[328]^u[31]^u[30]^u[25]^u[22]^u[17]^u[14]^u[12]^u[11]^u[4]^u[3]^u[1];
	y[160] = x[128]^x[299]^x[300]^x[305]^x[308]^x[313]^x[316]^x[318]^x[319]^x[326]^x[327]^x[329]^u[30]^u[29]^u[24]^u[21]^u[16]^u[13]^u[11]^u[10]^u[3]^u[2]^u[0];
	y[161] = x[129]^x[298]^x[299]^x[302]^x[304]^x[307]^x[309]^x[310]^x[314]^x[316]^x[317]^x[318]^x[323]^x[324]^x[325]^x[326]^x[328]^u[31]^u[30]^u[27]^u[25]^u[22]^u[20]^u[19]^u[15]^u[13]^u[12]^u[11]^u[6]^u[5]^u[4]^u[3]^u[1];
	y[162] = x[130]^x[298]^x[301]^x[302]^x[303]^x[304]^x[305]^x[306]^x[307]^x[308]^x[311]^x[315]^x[316]^x[317]^x[320]^x[323]^x[329]^u[31]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[18]^u[14]^u[13]^u[12]^u[9]^u[6]^u[0];
	y[163] = x[131]^x[298]^x[300]^x[301]^x[303]^x[305]^x[308]^x[309]^x[310]^x[312]^x[317]^x[319]^x[320]^x[321]^x[323]^x[325]^x[326]^x[327]^u[31]^u[29]^u[28]^u[26]^u[24]^u[21]^u[20]^u[19]^u[17]^u[12]^u[10]^u[9]^u[8]^u[6]^u[4]^u[3]^u[2];
	y[164] = x[132]^x[299]^x[301]^x[302]^x[304]^x[306]^x[309]^x[310]^x[311]^x[313]^x[318]^x[320]^x[321]^x[322]^x[324]^x[326]^x[327]^x[328]^u[30]^u[28]^u[27]^u[25]^u[23]^u[20]^u[19]^u[18]^u[16]^u[11]^u[9]^u[8]^u[7]^u[5]^u[3]^u[2]^u[1];
	y[165] = x[133]^x[298]^x[299]^x[301]^x[303]^x[304]^x[305]^x[306]^x[311]^x[312]^x[314]^x[316]^x[318]^x[320]^x[321]^x[322]^x[324]^x[326]^x[328]^x[329]^u[31]^u[30]^u[28]^u[26]^u[25]^u[24]^u[23]^u[18]^u[17]^u[15]^u[13]^u[11]^u[9]^u[8]^u[7]^u[5]^u[3]^u[1]^u[0];
	y[166] = x[134]^x[298]^x[301]^x[305]^x[310]^x[312]^x[313]^x[315]^x[316]^x[317]^x[318]^x[320]^x[321]^x[322]^x[324]^x[326]^x[329]^u[31]^u[28]^u[24]^u[19]^u[17]^u[16]^u[14]^u[13]^u[12]^u[11]^u[9]^u[8]^u[7]^u[5]^u[3]^u[0];
	y[167] = x[135]^x[299]^x[302]^x[306]^x[311]^x[313]^x[314]^x[316]^x[317]^x[318]^x[319]^x[321]^x[322]^x[323]^x[325]^x[327]^u[30]^u[27]^u[23]^u[18]^u[16]^u[15]^u[13]^u[12]^u[11]^u[10]^u[8]^u[7]^u[6]^u[4]^u[2];
	y[168] = x[136]^x[300]^x[303]^x[307]^x[312]^x[314]^x[315]^x[317]^x[318]^x[319]^x[320]^x[322]^x[323]^x[324]^x[326]^x[328]^u[29]^u[26]^u[22]^u[17]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[7]^u[6]^u[5]^u[3]^u[1];
	y[169] = x[137]^x[301]^x[304]^x[308]^x[313]^x[315]^x[316]^x[318]^x[319]^x[320]^x[321]^x[323]^x[324]^x[325]^x[327]^x[329]^u[28]^u[25]^u[21]^u[16]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4]^u[2]^u[0];
	y[170] = x[138]^x[302]^x[305]^x[309]^x[314]^x[316]^x[317]^x[319]^x[320]^x[321]^x[322]^x[324]^x[325]^x[326]^x[328]^u[27]^u[24]^u[20]^u[15]^u[13]^u[12]^u[10]^u[9]^u[8]^u[7]^u[5]^u[4]^u[3]^u[1];
	y[171] = x[139]^x[298]^x[299]^x[300]^x[301]^x[302]^x[303]^x[304]^x[307]^x[315]^x[316]^x[317]^x[319]^x[321]^x[322]^x[324]^x[329]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[22]^u[14]^u[13]^u[12]^u[10]^u[8]^u[7]^u[5]^u[0];
	y[172] = x[140]^x[298]^x[303]^x[305]^x[306]^x[307]^x[308]^x[310]^x[317]^x[319]^x[322]^x[324]^x[326]^x[327]^u[31]^u[26]^u[24]^u[23]^u[22]^u[21]^u[19]^u[12]^u[10]^u[7]^u[5]^u[3]^u[2];
	y[173] = x[141]^x[299]^x[304]^x[306]^x[307]^x[308]^x[309]^x[311]^x[318]^x[320]^x[323]^x[325]^x[327]^x[328]^u[30]^u[25]^u[23]^u[22]^u[21]^u[20]^u[18]^u[11]^u[9]^u[6]^u[4]^u[2]^u[1];
	y[174] = x[142]^x[298]^x[299]^x[301]^x[302]^x[304]^x[305]^x[306]^x[308]^x[309]^x[312]^x[316]^x[318]^x[320]^x[321]^x[323]^x[325]^x[327]^x[328]^x[329]^u[31]^u[30]^u[28]^u[27]^u[25]^u[24]^u[23]^u[21]^u[20]^u[17]^u[13]^u[11]^u[9]^u[8]^u[6]^u[4]^u[2]^u[1]^u[0];
	y[175] = x[143]^x[299]^x[300]^x[302]^x[303]^x[305]^x[306]^x[307]^x[309]^x[310]^x[313]^x[317]^x[319]^x[321]^x[322]^x[324]^x[326]^x[328]^x[329]^u[30]^u[29]^u[27]^u[26]^u[24]^u[23]^u[22]^u[20]^u[19]^u[16]^u[12]^u[10]^u[8]^u[7]^u[5]^u[3]^u[1]^u[0];
	y[176] = x[144]^x[300]^x[301]^x[303]^x[304]^x[306]^x[307]^x[308]^x[310]^x[311]^x[314]^x[318]^x[320]^x[322]^x[323]^x[325]^x[327]^x[329]^u[29]^u[28]^u[26]^u[25]^u[23]^u[22]^u[21]^u[19]^u[18]^u[15]^u[11]^u[9]^u[7]^u[6]^u[4]^u[2]^u[0];
	y[177] = x[145]^x[301]^x[302]^x[304]^x[305]^x[307]^x[308]^x[309]^x[311]^x[312]^x[315]^x[319]^x[321]^x[323]^x[324]^x[326]^x[328]^u[28]^u[27]^u[25]^u[24]^u[22]^u[21]^u[20]^u[18]^u[17]^u[14]^u[10]^u[8]^u[6]^u[5]^u[3]^u[1];
	y[178] = x[146]^x[298]^x[299]^x[300]^x[301]^x[303]^x[304]^x[305]^x[307]^x[308]^x[309]^x[312]^x[313]^x[318]^x[319]^x[322]^x[323]^x[326]^x[329]^u[31]^u[30]^u[29]^u[28]^u[26]^u[25]^u[24]^u[22]^u[21]^u[20]^u[17]^u[16]^u[11]^u[10]^u[7]^u[6]^u[3]^u[0];
	y[179] = x[147]^x[298]^x[305]^x[307]^x[308]^x[309]^x[313]^x[314]^x[316]^x[318]^x[325]^x[326]^u[31]^u[24]^u[22]^u[21]^u[20]^u[16]^u[15]^u[13]^u[11]^u[4]^u[3];
	y[180] = x[148]^x[299]^x[306]^x[308]^x[309]^x[310]^x[314]^x[315]^x[317]^x[319]^x[326]^x[327]^u[30]^u[23]^u[21]^u[20]^u[19]^u[15]^u[14]^u[12]^u[10]^u[3]^u[2];
	y[181] = x[149]^x[300]^x[307]^x[309]^x[310]^x[311]^x[315]^x[316]^x[318]^x[320]^x[327]^x[328]^u[29]^u[22]^u[20]^u[19]^u[18]^u[14]^u[13]^u[11]^u[9]^u[2]^u[1];
	y[182] = x[150]^x[301]^x[308]^x[310]^x[311]^x[312]^x[316]^x[317]^x[319]^x[321]^x[328]^x[329]^u[28]^u[21]^u[19]^u[18]^u[17]^u[13]^u[12]^u[10]^u[8]^u[1]^u[0];
	y[183] = x[151]^x[302]^x[309]^x[311]^x[312]^x[313]^x[317]^x[318]^x[320]^x[322]^x[329]^u[27]^u[20]^u[18]^u[17]^u[16]^u[12]^u[11]^u[9]^u[7]^u[0];
	y[184] = x[152]^x[298]^x[299]^x[300]^x[301]^x[302]^x[303]^x[304]^x[306]^x[307]^x[312]^x[313]^x[314]^x[316]^x[320]^x[321]^x[324]^x[325]^x[326]^x[327]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[23]^u[22]^u[17]^u[16]^u[15]^u[13]^u[9]^u[8]^u[5]^u[4]^u[3]^u[2];
	y[185] = x[153]^x[298]^x[303]^x[305]^x[306]^x[308]^x[310]^x[313]^x[314]^x[315]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[328]^u[31]^u[26]^u[24]^u[23]^u[21]^u[19]^u[16]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[1];
	y[186] = x[154]^x[299]^x[304]^x[306]^x[307]^x[309]^x[311]^x[314]^x[315]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[325]^x[329]^u[30]^u[25]^u[23]^u[22]^u[20]^u[18]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[0];
	y[187] = x[155]^x[298]^x[299]^x[301]^x[302]^x[304]^x[305]^x[306]^x[308]^x[312]^x[315]^x[317]^x[321]^x[322]^x[327]^u[31]^u[30]^u[28]^u[27]^u[25]^u[24]^u[23]^u[21]^u[17]^u[14]^u[12]^u[8]^u[7]^u[2];
	y[188] = x[156]^x[299]^x[300]^x[302]^x[303]^x[305]^x[306]^x[307]^x[309]^x[313]^x[316]^x[318]^x[322]^x[323]^x[328]^u[30]^u[29]^u[27]^u[26]^u[24]^u[23]^u[22]^u[20]^u[16]^u[13]^u[11]^u[7]^u[6]^u[1];
	y[189] = x[157]^x[298]^x[299]^x[302]^x[303]^x[308]^x[314]^x[316]^x[317]^x[318]^x[320]^x[325]^x[326]^x[327]^x[329]^u[31]^u[30]^u[27]^u[26]^u[21]^u[15]^u[13]^u[12]^u[11]^u[9]^u[4]^u[3]^u[2]^u[0];
	y[190] = x[158]^x[299]^x[300]^x[303]^x[304]^x[309]^x[315]^x[317]^x[318]^x[319]^x[321]^x[326]^x[327]^x[328]^u[30]^u[29]^u[26]^u[25]^u[20]^u[14]^u[12]^u[11]^u[10]^u[8]^u[3]^u[2]^u[1];
	y[191] = x[159]^x[300]^x[301]^x[304]^x[305]^x[310]^x[316]^x[318]^x[319]^x[320]^x[322]^x[327]^x[328]^x[329]^u[29]^u[28]^u[25]^u[24]^u[19]^u[13]^u[11]^u[10]^u[9]^u[7]^u[2]^u[1]^u[0];
	y[192] = x[160]^x[298]^x[299]^x[300]^x[304]^x[305]^x[307]^x[310]^x[311]^x[316]^x[317]^x[318]^x[321]^x[324]^x[325]^x[326]^x[327]^x[328]^x[329]^u[31]^u[30]^u[29]^u[25]^u[24]^u[22]^u[19]^u[18]^u[13]^u[12]^u[11]^u[8]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[193] = x[161]^x[298]^x[302]^x[304]^x[305]^x[307]^x[308]^x[310]^x[311]^x[312]^x[316]^x[317]^x[320]^x[322]^x[323]^x[324]^x[328]^x[329]^u[31]^u[27]^u[25]^u[24]^u[22]^u[21]^u[19]^u[18]^u[17]^u[13]^u[12]^u[9]^u[7]^u[6]^u[5]^u[1]^u[0];
	y[194] = x[162]^x[299]^x[303]^x[305]^x[306]^x[308]^x[309]^x[311]^x[312]^x[313]^x[317]^x[318]^x[321]^x[323]^x[324]^x[325]^x[329]^u[30]^u[26]^u[24]^u[23]^u[21]^u[20]^u[18]^u[17]^u[16]^u[12]^u[11]^u[8]^u[6]^u[5]^u[4]^u[0];
	y[195] = x[163]^x[298]^x[299]^x[301]^x[302]^x[309]^x[312]^x[313]^x[314]^x[316]^x[320]^x[322]^x[323]^x[327]^u[31]^u[30]^u[28]^u[27]^u[20]^u[17]^u[16]^u[15]^u[13]^u[9]^u[7]^u[6]^u[2];
	y[196] = x[164]^x[298]^x[301]^x[303]^x[304]^x[306]^x[307]^x[313]^x[314]^x[315]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[325]^x[326]^x[327]^x[328]^u[31]^u[28]^u[26]^u[25]^u[23]^u[22]^u[16]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[4]^u[3]^u[2]^u[1];
	y[197] = x[165]^x[299]^x[302]^x[304]^x[305]^x[307]^x[308]^x[314]^x[315]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[326]^x[327]^x[328]^x[329]^u[30]^u[27]^u[25]^u[24]^u[22]^u[21]^u[15]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[3]^u[2]^u[1]^u[0];
	y[198] = x[166]^x[300]^x[303]^x[305]^x[306]^x[308]^x[309]^x[315]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[327]^x[328]^x[329]^u[29]^u[26]^u[24]^u[23]^u[21]^u[20]^u[14]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[2]^u[1]^u[0];
	y[199] = x[167]^x[301]^x[304]^x[306]^x[307]^x[309]^x[310]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[328]^x[329]^u[28]^u[25]^u[23]^u[22]^u[20]^u[19]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[1]^u[0];
	y[200] = x[168]^x[298]^x[299]^x[300]^x[301]^x[304]^x[305]^x[306]^x[308]^x[311]^x[316]^x[317]^x[321]^x[322]^x[326]^x[327]^x[329]^u[31]^u[30]^u[29]^u[28]^u[25]^u[24]^u[23]^u[21]^u[18]^u[13]^u[12]^u[8]^u[7]^u[3]^u[2]^u[0];
	y[201] = x[169]^x[299]^x[300]^x[301]^x[302]^x[305]^x[306]^x[307]^x[309]^x[312]^x[317]^x[318]^x[322]^x[323]^x[327]^x[328]^u[30]^u[29]^u[28]^u[27]^u[24]^u[23]^u[22]^u[20]^u[17]^u[12]^u[11]^u[7]^u[6]^u[2]^u[1];
	y[202] = x[170]^x[298]^x[299]^x[303]^x[304]^x[308]^x[313]^x[316]^x[320]^x[325]^x[326]^x[327]^x[328]^x[329]^u[31]^u[30]^u[26]^u[25]^u[21]^u[16]^u[13]^u[9]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[203] = x[171]^x[298]^x[301]^x[302]^x[305]^x[306]^x[307]^x[309]^x[310]^x[314]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[323]^x[324]^x[325]^x[328]^x[329]^u[31]^u[28]^u[27]^u[24]^u[23]^u[22]^u[20]^u[19]^u[15]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4]^u[1]^u[0];
	y[204] = x[172]^x[298]^x[300]^x[301]^x[303]^x[304]^x[308]^x[311]^x[315]^x[316]^x[317]^x[321]^x[322]^x[323]^x[327]^x[329]^u[31]^u[29]^u[28]^u[26]^u[25]^u[21]^u[18]^u[14]^u[13]^u[12]^u[8]^u[7]^u[6]^u[2]^u[0];
	y[205] = x[173]^x[298]^x[300]^x[305]^x[306]^x[307]^x[309]^x[310]^x[312]^x[317]^x[319]^x[320]^x[322]^x[325]^x[326]^x[327]^x[328]^u[31]^u[29]^u[24]^u[23]^u[22]^u[20]^u[19]^u[17]^u[12]^u[10]^u[9]^u[7]^u[4]^u[3]^u[2]^u[1];
	y[206] = x[174]^x[299]^x[301]^x[306]^x[307]^x[308]^x[310]^x[311]^x[313]^x[318]^x[320]^x[321]^x[323]^x[326]^x[327]^x[328]^x[329]^u[30]^u[28]^u[23]^u[22]^u[21]^u[19]^u[18]^u[16]^u[11]^u[9]^u[8]^u[6]^u[3]^u[2]^u[1]^u[0];
	y[207] = x[175]^x[300]^x[302]^x[307]^x[308]^x[309]^x[311]^x[312]^x[314]^x[319]^x[321]^x[322]^x[324]^x[327]^x[328]^x[329]^u[29]^u[27]^u[22]^u[21]^u[20]^u[18]^u[17]^u[15]^u[10]^u[8]^u[7]^u[5]^u[2]^u[1]^u[0];
	y[208] = x[176]^x[298]^x[299]^x[300]^x[302]^x[303]^x[304]^x[306]^x[307]^x[308]^x[309]^x[312]^x[313]^x[315]^x[316]^x[318]^x[319]^x[322]^x[324]^x[326]^x[327]^x[328]^x[329]^u[31]^u[30]^u[29]^u[27]^u[26]^u[25]^u[23]^u[22]^u[21]^u[20]^u[17]^u[16]^u[14]^u[13]^u[11]^u[10]^u[7]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[209] = x[177]^x[299]^x[300]^x[301]^x[303]^x[304]^x[305]^x[307]^x[308]^x[309]^x[310]^x[313]^x[314]^x[316]^x[317]^x[319]^x[320]^x[323]^x[325]^x[327]^x[328]^x[329]^u[30]^u[29]^u[28]^u[26]^u[25]^u[24]^u[22]^u[21]^u[20]^u[19]^u[16]^u[15]^u[13]^u[12]^u[10]^u[9]^u[6]^u[4]^u[2]^u[1]^u[0];
	y[210] = x[178]^x[298]^x[299]^x[305]^x[307]^x[308]^x[309]^x[311]^x[314]^x[315]^x[316]^x[317]^x[319]^x[321]^x[323]^x[325]^x[327]^x[328]^x[329]^u[31]^u[30]^u[24]^u[22]^u[21]^u[20]^u[18]^u[15]^u[14]^u[13]^u[12]^u[10]^u[8]^u[6]^u[4]^u[2]^u[1]^u[0];
	y[211] = x[179]^x[298]^x[301]^x[302]^x[304]^x[307]^x[308]^x[309]^x[312]^x[315]^x[317]^x[319]^x[322]^x[323]^x[325]^x[327]^x[328]^x[329]^u[31]^u[28]^u[27]^u[25]^u[22]^u[21]^u[20]^u[17]^u[14]^u[12]^u[10]^u[7]^u[6]^u[4]^u[2]^u[1]^u[0];
	y[212] = x[180]^x[299]^x[302]^x[303]^x[305]^x[308]^x[309]^x[310]^x[313]^x[316]^x[318]^x[320]^x[323]^x[324]^x[326]^x[328]^x[329]^u[30]^u[27]^u[26]^u[24]^u[21]^u[20]^u[19]^u[16]^u[13]^u[11]^u[9]^u[6]^u[5]^u[3]^u[1]^u[0];
	y[213] = x[181]^x[300]^x[303]^x[304]^x[306]^x[309]^x[310]^x[311]^x[314]^x[317]^x[319]^x[321]^x[324]^x[325]^x[327]^x[329]^u[29]^u[26]^u[25]^u[23]^u[20]^u[19]^u[18]^u[15]^u[12]^u[10]^u[8]^u[5]^u[4]^u[2]^u[0];
	y[214] = x[182]^x[298]^x[299]^x[300]^x[302]^x[305]^x[306]^x[311]^x[312]^x[315]^x[316]^x[319]^x[322]^x[323]^x[324]^x[327]^x[328]^u[31]^u[30]^u[29]^u[27]^u[24]^u[23]^u[18]^u[17]^u[14]^u[13]^u[10]^u[7]^u[6]^u[5]^u[2]^u[1];
	y[215] = x[183]^x[299]^x[300]^x[301]^x[303]^x[306]^x[307]^x[312]^x[313]^x[316]^x[317]^x[320]^x[323]^x[324]^x[325]^x[328]^x[329]^u[30]^u[29]^u[28]^u[26]^u[23]^u[22]^u[17]^u[16]^u[13]^u[12]^u[9]^u[6]^u[5]^u[4]^u[1]^u[0];
	y[216] = x[184]^x[300]^x[301]^x[302]^x[304]^x[307]^x[308]^x[313]^x[314]^x[317]^x[318]^x[321]^x[324]^x[325]^x[326]^x[329]^u[29]^u[28]^u[27]^u[25]^u[22]^u[21]^u[16]^u[15]^u[12]^u[11]^u[8]^u[5]^u[4]^u[3]^u[0];
	y[217] = x[185]^x[301]^x[302]^x[303]^x[305]^x[308]^x[309]^x[314]^x[315]^x[318]^x[319]^x[322]^x[325]^x[326]^x[327]^u[28]^u[27]^u[26]^u[24]^u[21]^u[20]^u[15]^u[14]^u[11]^u[10]^u[7]^u[4]^u[3]^u[2];
	y[218] = x[186]^x[298]^x[299]^x[300]^x[301]^x[303]^x[307]^x[309]^x[315]^x[318]^x[324]^x[325]^x[328]^u[31]^u[30]^u[29]^u[28]^u[26]^u[22]^u[20]^u[14]^u[11]^u[5]^u[4]^u[1];
	y[219] = x[187]^x[298]^x[306]^x[307]^x[308]^x[318]^x[320]^x[323]^x[324]^x[327]^x[329]^u[31]^u[23]^u[22]^u[21]^u[11]^u[9]^u[6]^u[5]^u[2]^u[0];
	y[220] = x[188]^x[299]^x[307]^x[308]^x[309]^x[319]^x[321]^x[324]^x[325]^x[328]^u[30]^u[22]^u[21]^u[20]^u[10]^u[8]^u[5]^u[4]^u[1];
	y[221] = x[189]^x[300]^x[308]^x[309]^x[310]^x[320]^x[322]^x[325]^x[326]^x[329]^u[29]^u[21]^u[20]^u[19]^u[9]^u[7]^u[4]^u[3]^u[0];
	y[222] = x[190]^x[301]^x[309]^x[310]^x[311]^x[321]^x[323]^x[326]^x[327]^u[28]^u[20]^u[19]^u[18]^u[8]^u[6]^u[3]^u[2];
	y[223] = x[191]^x[298]^x[299]^x[300]^x[301]^x[304]^x[306]^x[307]^x[311]^x[312]^x[316]^x[318]^x[319]^x[320]^x[322]^x[323]^x[325]^x[326]^x[328]^u[31]^u[30]^u[29]^u[28]^u[25]^u[23]^u[22]^u[18]^u[17]^u[13]^u[11]^u[10]^u[9]^u[7]^u[6]^u[4]^u[3]^u[1];
	y[224] = x[192]^x[298]^x[304]^x[305]^x[306]^x[308]^x[310]^x[312]^x[313]^x[316]^x[317]^x[318]^x[321]^x[325]^x[329]^u[31]^u[25]^u[24]^u[23]^u[21]^u[19]^u[17]^u[16]^u[13]^u[12]^u[11]^u[8]^u[4]^u[0];
	y[225] = x[193]^x[299]^x[305]^x[306]^x[307]^x[309]^x[311]^x[313]^x[314]^x[317]^x[318]^x[319]^x[322]^x[326]^u[30]^u[24]^u[23]^u[22]^u[20]^u[18]^u[16]^u[15]^u[12]^u[11]^u[10]^u[7]^u[3];
	y[226] = x[194]^x[300]^x[306]^x[307]^x[308]^x[310]^x[312]^x[314]^x[315]^x[318]^x[319]^x[320]^x[323]^x[327]^u[29]^u[23]^u[22]^u[21]^u[19]^u[17]^u[15]^u[14]^u[11]^u[10]^u[9]^u[6]^u[2];
	y[227] = x[195]^x[301]^x[307]^x[308]^x[309]^x[311]^x[313]^x[315]^x[316]^x[319]^x[320]^x[321]^x[324]^x[328]^u[28]^u[22]^u[21]^u[20]^u[18]^u[16]^u[14]^u[13]^u[10]^u[9]^u[8]^u[5]^u[1];
	y[228] = x[196]^x[298]^x[299]^x[300]^x[301]^x[304]^x[306]^x[307]^x[308]^x[309]^x[312]^x[314]^x[317]^x[318]^x[319]^x[321]^x[322]^x[323]^x[324]^x[326]^x[327]^x[329]^u[31]^u[30]^u[29]^u[28]^u[25]^u[23]^u[22]^u[21]^u[20]^u[17]^u[15]^u[12]^u[11]^u[10]^u[8]^u[7]^u[6]^u[5]^u[3]^u[2]^u[0];
	y[229] = x[197]^x[299]^x[300]^x[301]^x[302]^x[305]^x[307]^x[308]^x[309]^x[310]^x[313]^x[315]^x[318]^x[319]^x[320]^x[322]^x[323]^x[324]^x[325]^x[327]^x[328]^u[30]^u[29]^u[28]^u[27]^u[24]^u[22]^u[21]^u[20]^u[19]^u[16]^u[14]^u[11]^u[10]^u[9]^u[7]^u[6]^u[5]^u[4]^u[2]^u[1];
	y[230] = x[198]^x[300]^x[301]^x[302]^x[303]^x[306]^x[308]^x[309]^x[310]^x[311]^x[314]^x[316]^x[319]^x[320]^x[321]^x[323]^x[324]^x[325]^x[326]^x[328]^x[329]^u[29]^u[28]^u[27]^u[26]^u[23]^u[21]^u[20]^u[19]^u[18]^u[15]^u[13]^u[10]^u[9]^u[8]^u[6]^u[5]^u[4]^u[3]^u[1]^u[0];
	y[231] = x[199]^x[301]^x[302]^x[303]^x[304]^x[307]^x[309]^x[310]^x[311]^x[312]^x[315]^x[317]^x[320]^x[321]^x[322]^x[324]^x[325]^x[326]^x[327]^x[329]^u[28]^u[27]^u[26]^u[25]^u[22]^u[20]^u[19]^u[18]^u[17]^u[14]^u[12]^u[9]^u[8]^u[7]^u[5]^u[4]^u[3]^u[2]^u[0];
	y[232] = x[200]^x[302]^x[303]^x[304]^x[305]^x[308]^x[310]^x[311]^x[312]^x[313]^x[316]^x[318]^x[321]^x[322]^x[323]^x[325]^x[326]^x[327]^x[328]^u[27]^u[26]^u[25]^u[24]^u[21]^u[19]^u[18]^u[17]^u[16]^u[13]^u[11]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1];
	y[233] = x[201]^x[303]^x[304]^x[305]^x[306]^x[309]^x[311]^x[312]^x[313]^x[314]^x[317]^x[319]^x[322]^x[323]^x[324]^x[326]^x[327]^x[328]^x[329]^u[26]^u[25]^u[24]^u[23]^u[20]^u[18]^u[17]^u[16]^u[15]^u[12]^u[10]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1]^u[0];
	y[234] = x[202]^x[298]^x[299]^x[300]^x[301]^x[302]^x[305]^x[312]^x[313]^x[314]^x[315]^x[316]^x[319]^x[326]^x[328]^x[329]^u[31]^u[30]^u[29]^u[28]^u[27]^u[24]^u[17]^u[16]^u[15]^u[14]^u[13]^u[10]^u[3]^u[1]^u[0];
	y[235] = x[203]^x[299]^x[300]^x[301]^x[302]^x[303]^x[306]^x[313]^x[314]^x[315]^x[316]^x[317]^x[320]^x[327]^x[329]^u[30]^u[29]^u[28]^u[27]^u[26]^u[23]^u[16]^u[15]^u[14]^u[13]^u[12]^u[9]^u[2]^u[0];
	y[236] = x[204]^x[300]^x[301]^x[302]^x[303]^x[304]^x[307]^x[314]^x[315]^x[316]^x[317]^x[318]^x[321]^x[328]^u[29]^u[28]^u[27]^u[26]^u[25]^u[22]^u[15]^u[14]^u[13]^u[12]^u[11]^u[8]^u[1];
	y[237] = x[205]^x[298]^x[299]^x[300]^x[303]^x[305]^x[306]^x[307]^x[308]^x[310]^x[315]^x[317]^x[320]^x[322]^x[323]^x[324]^x[325]^x[326]^x[327]^x[329]^u[31]^u[30]^u[29]^u[26]^u[24]^u[23]^u[22]^u[21]^u[19]^u[14]^u[12]^u[9]^u[7]^u[6]^u[5]^u[4]^u[3]^u[2]^u[0];
	y[238] = x[206]^x[299]^x[300]^x[301]^x[304]^x[306]^x[307]^x[308]^x[309]^x[311]^x[316]^x[318]^x[321]^x[323]^x[324]^x[325]^x[326]^x[327]^x[328]^u[30]^u[29]^u[28]^u[25]^u[23]^u[22]^u[21]^u[20]^u[18]^u[13]^u[11]^u[8]^u[6]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[239] = x[207]^x[300]^x[301]^x[302]^x[305]^x[307]^x[308]^x[309]^x[310]^x[312]^x[317]^x[319]^x[322]^x[324]^x[325]^x[326]^x[327]^x[328]^x[329]^u[29]^u[28]^u[27]^u[24]^u[22]^u[21]^u[20]^u[19]^u[17]^u[12]^u[10]^u[7]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[240] = x[208]^x[301]^x[302]^x[303]^x[306]^x[308]^x[309]^x[310]^x[311]^x[313]^x[318]^x[320]^x[323]^x[325]^x[326]^x[327]^x[328]^x[329]^u[28]^u[27]^u[26]^u[23]^u[21]^u[20]^u[19]^u[18]^u[16]^u[11]^u[9]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[241] = x[209]^x[298]^x[299]^x[300]^x[301]^x[303]^x[306]^x[309]^x[311]^x[312]^x[314]^x[316]^x[318]^x[320]^x[321]^x[323]^x[325]^x[328]^x[329]^u[31]^u[30]^u[29]^u[28]^u[26]^u[23]^u[20]^u[18]^u[17]^u[15]^u[13]^u[11]^u[9]^u[8]^u[6]^u[4]^u[1]^u[0];
	y[242] = x[210]^x[299]^x[300]^x[301]^x[302]^x[304]^x[307]^x[310]^x[312]^x[313]^x[315]^x[317]^x[319]^x[321]^x[322]^x[324]^x[326]^x[329]^u[30]^u[29]^u[28]^u[27]^u[25]^u[22]^u[19]^u[17]^u[16]^u[14]^u[12]^u[10]^u[8]^u[7]^u[5]^u[3]^u[0];
	y[243] = x[211]^x[300]^x[301]^x[302]^x[303]^x[305]^x[308]^x[311]^x[313]^x[314]^x[316]^x[318]^x[320]^x[322]^x[323]^x[325]^x[327]^u[29]^u[28]^u[27]^u[26]^u[24]^u[21]^u[18]^u[16]^u[15]^u[13]^u[11]^u[9]^u[7]^u[6]^u[4]^u[2];
	y[244] = x[212]^x[301]^x[302]^x[303]^x[304]^x[306]^x[309]^x[312]^x[314]^x[315]^x[317]^x[319]^x[321]^x[323]^x[324]^x[326]^x[328]^u[28]^u[27]^u[26]^u[25]^u[23]^u[20]^u[17]^u[15]^u[14]^u[12]^u[10]^u[8]^u[6]^u[5]^u[3]^u[1];
	y[245] = x[213]^x[298]^x[299]^x[300]^x[301]^x[303]^x[305]^x[306]^x[313]^x[315]^x[319]^x[322]^x[323]^x[326]^x[329]^u[31]^u[30]^u[29]^u[28]^u[26]^u[24]^u[23]^u[16]^u[14]^u[10]^u[7]^u[6]^u[3]^u[0];
	y[246] = x[214]^x[299]^x[300]^x[301]^x[302]^x[304]^x[306]^x[307]^x[314]^x[316]^x[320]^x[323]^x[324]^x[327]^u[30]^u[29]^u[28]^u[27]^u[25]^u[23]^u[22]^u[15]^u[13]^u[9]^u[6]^u[5]^u[2];
	y[247] = x[215]^x[300]^x[301]^x[302]^x[303]^x[305]^x[307]^x[308]^x[315]^x[317]^x[321]^x[324]^x[325]^x[328]^u[29]^u[28]^u[27]^u[26]^u[24]^u[22]^u[21]^u[14]^u[12]^u[8]^u[5]^u[4]^u[1];
	y[248] = x[216]^x[301]^x[302]^x[303]^x[304]^x[306]^x[308]^x[309]^x[316]^x[318]^x[322]^x[325]^x[326]^x[329]^u[28]^u[27]^u[26]^u[25]^u[23]^u[21]^u[20]^u[13]^u[11]^u[7]^u[4]^u[3]^u[0];
	y[249] = x[217]^x[298]^x[299]^x[300]^x[301]^x[303]^x[305]^x[306]^x[309]^x[316]^x[317]^x[318]^x[320]^x[324]^x[325]^u[31]^u[30]^u[29]^u[28]^u[26]^u[24]^u[23]^u[20]^u[13]^u[12]^u[11]^u[9]^u[5]^u[4];
	y[250] = x[218]^x[298]^x[316]^x[317]^x[320]^x[321]^x[323]^x[324]^x[327]^u[31]^u[13]^u[12]^u[9]^u[8]^u[6]^u[5]^u[2];
	y[251] = x[219]^x[299]^x[317]^x[318]^x[321]^x[322]^x[324]^x[325]^x[328]^u[30]^u[12]^u[11]^u[8]^u[7]^u[5]^u[4]^u[1];
	y[252] = x[220]^x[300]^x[318]^x[319]^x[322]^x[323]^x[325]^x[326]^x[329]^u[29]^u[11]^u[10]^u[7]^u[6]^u[4]^u[3]^u[0];
	y[253] = x[221]^x[301]^x[319]^x[320]^x[323]^x[324]^x[326]^x[327]^u[28]^u[10]^u[9]^u[6]^u[5]^u[3]^u[2];
	y[254] = x[222]^x[298]^x[299]^x[300]^x[301]^x[304]^x[306]^x[307]^x[310]^x[316]^x[318]^x[319]^x[321]^x[323]^x[326]^x[328]^u[31]^u[30]^u[29]^u[28]^u[25]^u[23]^u[22]^u[19]^u[13]^u[11]^u[10]^u[8]^u[6]^u[3]^u[1];
	y[255] = x[223]^x[299]^x[300]^x[301]^x[302]^x[305]^x[307]^x[308]^x[311]^x[317]^x[319]^x[320]^x[322]^x[324]^x[327]^x[329]^u[30]^u[29]^u[28]^u[27]^u[24]^u[22]^u[21]^u[18]^u[12]^u[10]^u[9]^u[7]^u[5]^u[2]^u[0];
	y[256] = x[224]^x[300]^x[301]^x[302]^x[303]^x[306]^x[308]^x[309]^x[312]^x[318]^x[320]^x[321]^x[323]^x[325]^x[328]^u[29]^u[28]^u[27]^u[26]^u[23]^u[21]^u[20]^u[17]^u[11]^u[9]^u[8]^u[6]^u[4]^u[1];
	y[257] = x[225]^x[301]^x[302]^x[303]^x[304]^x[307]^x[309]^x[310]^x[313]^x[319]^x[321]^x[322]^x[324]^x[326]^x[329]^u[28]^u[27]^u[26]^u[25]^u[22]^u[20]^u[19]^u[16]^u[10]^u[8]^u[7]^u[5]^u[3]^u[0];
	y[258] = x[226]^x[298]^x[299]^x[300]^x[301]^x[303]^x[305]^x[306]^x[307]^x[308]^x[311]^x[314]^x[316]^x[318]^x[319]^x[322]^x[324]^x[326]^u[31]^u[30]^u[29]^u[28]^u[26]^u[24]^u[23]^u[22]^u[21]^u[18]^u[15]^u[13]^u[11]^u[10]^u[7]^u[5]^u[3];
	y[259] = x[227]^x[298]^x[308]^x[309]^x[310]^x[312]^x[315]^x[316]^x[317]^x[318]^x[324]^x[326]^u[31]^u[21]^u[20]^u[19]^u[17]^u[14]^u[13]^u[12]^u[11]^u[5]^u[3];
	y[260] = x[228]^x[299]^x[309]^x[310]^x[311]^x[313]^x[316]^x[317]^x[318]^x[319]^x[325]^x[327]^u[30]^u[20]^u[19]^u[18]^u[16]^u[13]^u[12]^u[11]^u[10]^u[4]^u[2];
	y[261] = x[229]^x[300]^x[310]^x[311]^x[312]^x[314]^x[317]^x[318]^x[319]^x[320]^x[326]^x[328]^u[29]^u[19]^u[18]^u[17]^u[15]^u[12]^u[11]^u[10]^u[9]^u[3]^u[1];
	y[262] = x[230]^x[298]^x[299]^x[300]^x[302]^x[304]^x[306]^x[307]^x[310]^x[311]^x[312]^x[313]^x[315]^x[316]^x[321]^x[323]^x[324]^x[325]^x[326]^x[329]^u[31]^u[30]^u[29]^u[27]^u[25]^u[23]^u[22]^u[19]^u[18]^u[17]^u[16]^u[14]^u[13]^u[8]^u[6]^u[5]^u[4]^u[3]^u[0];
	y[263] = x[231]^x[299]^x[300]^x[301]^x[303]^x[305]^x[307]^x[308]^x[311]^x[312]^x[313]^x[314]^x[316]^x[317]^x[322]^x[324]^x[325]^x[326]^x[327]^u[30]^u[29]^u[28]^u[26]^u[24]^u[22]^u[21]^u[18]^u[17]^u[16]^u[15]^u[13]^u[12]^u[7]^u[5]^u[4]^u[3]^u[2];
	y[264] = x[232]^x[298]^x[299]^x[307]^x[308]^x[309]^x[310]^x[312]^x[313]^x[314]^x[315]^x[316]^x[317]^x[319]^x[320]^x[324]^x[328]^u[31]^u[30]^u[22]^u[21]^u[20]^u[19]^u[17]^u[16]^u[15]^u[14]^u[13]^u[12]^u[10]^u[9]^u[5]^u[1];
	y[265] = x[233]^x[298]^x[301]^x[302]^x[304]^x[306]^x[307]^x[308]^x[309]^x[311]^x[313]^x[314]^x[315]^x[317]^x[319]^x[321]^x[323]^x[324]^x[326]^x[327]^x[329]^u[31]^u[28]^u[27]^u[25]^u[23]^u[22]^u[21]^u[20]^u[18]^u[16]^u[15]^u[14]^u[12]^u[10]^u[8]^u[6]^u[5]^u[3]^u[2]^u[0];
	y[266] = x[234]^x[298]^x[300]^x[301]^x[303]^x[304]^x[305]^x[306]^x[308]^x[309]^x[312]^x[314]^x[315]^x[319]^x[322]^x[323]^x[326]^x[328]^u[31]^u[29]^u[28]^u[26]^u[25]^u[24]^u[23]^u[21]^u[20]^u[17]^u[15]^u[14]^u[10]^u[7]^u[6]^u[3]^u[1];
	y[267] = x[235]^x[298]^x[300]^x[305]^x[309]^x[313]^x[315]^x[318]^x[319]^x[325]^x[326]^x[329]^u[31]^u[29]^u[24]^u[20]^u[16]^u[14]^u[11]^u[10]^u[4]^u[3]^u[0];
	y[268] = x[236]^x[298]^x[300]^x[302]^x[304]^x[307]^x[314]^x[318]^x[323]^x[324]^x[325]^u[31]^u[29]^u[27]^u[25]^u[22]^u[15]^u[11]^u[6]^u[5]^u[4];
	y[269] = x[237]^x[298]^x[300]^x[302]^x[303]^x[304]^x[305]^x[306]^x[307]^x[308]^x[310]^x[315]^x[316]^x[318]^x[320]^x[323]^x[327]^u[31]^u[29]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[19]^u[14]^u[13]^u[11]^u[9]^u[6]^u[2];
	y[270] = x[238]^x[299]^x[301]^x[303]^x[304]^x[305]^x[306]^x[307]^x[308]^x[309]^x[311]^x[316]^x[317]^x[319]^x[321]^x[324]^x[328]^u[30]^u[28]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[20]^u[18]^u[13]^u[12]^u[10]^u[8]^u[5]^u[1];
	y[271] = x[239]^x[298]^x[299]^x[301]^x[305]^x[308]^x[309]^x[312]^x[316]^x[317]^x[319]^x[322]^x[323]^x[324]^x[326]^x[327]^x[329]^u[31]^u[30]^u[28]^u[24]^u[21]^u[20]^u[17]^u[13]^u[12]^u[10]^u[7]^u[6]^u[5]^u[3]^u[2]^u[0];
	y[272] = x[240]^x[298]^x[301]^x[304]^x[307]^x[309]^x[313]^x[316]^x[317]^x[319]^x[326]^x[328]^u[31]^u[28]^u[25]^u[22]^u[20]^u[16]^u[13]^u[12]^u[10]^u[3]^u[1];
	y[273] = x[241]^x[299]^x[302]^x[305]^x[308]^x[310]^x[314]^x[317]^x[318]^x[320]^x[327]^x[329]^u[30]^u[27]^u[24]^u[21]^u[19]^u[15]^u[12]^u[11]^u[9]^u[2]^u[0];
	y[274] = x[242]^x[300]^x[303]^x[306]^x[309]^x[311]^x[315]^x[318]^x[319]^x[321]^x[328]^u[29]^u[26]^u[23]^u[20]^u[18]^u[14]^u[11]^u[10]^u[8]^u[1];
	y[275] = x[243]^x[301]^x[304]^x[307]^x[310]^x[312]^x[316]^x[319]^x[320]^x[322]^x[329]^u[28]^u[25]^u[22]^u[19]^u[17]^u[13]^u[10]^u[9]^u[7]^u[0];
	y[276] = x[244]^x[302]^x[305]^x[308]^x[311]^x[313]^x[317]^x[320]^x[321]^x[323]^u[27]^u[24]^u[21]^u[18]^u[16]^u[12]^u[9]^u[8]^u[6];
	y[277] = x[245]^x[298]^x[299]^x[300]^x[301]^x[302]^x[303]^x[304]^x[307]^x[309]^x[310]^x[312]^x[314]^x[316]^x[319]^x[320]^x[321]^x[322]^x[323]^x[325]^x[326]^x[327]^u[31]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[22]^u[20]^u[19]^u[17]^u[15]^u[13]^u[10]^u[9]^u[8]^u[7]^u[6]^u[4]^u[3]^u[2];
	y[278] = x[246]^x[299]^x[300]^x[301]^x[302]^x[303]^x[304]^x[305]^x[308]^x[310]^x[311]^x[313]^x[315]^x[317]^x[320]^x[321]^x[322]^x[323]^x[324]^x[326]^x[327]^x[328]^u[30]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[21]^u[19]^u[18]^u[16]^u[14]^u[12]^u[9]^u[8]^u[7]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[279] = x[247]^x[300]^x[301]^x[302]^x[303]^x[304]^x[305]^x[306]^x[309]^x[311]^x[312]^x[314]^x[316]^x[318]^x[321]^x[322]^x[323]^x[324]^x[325]^x[327]^x[328]^x[329]^u[29]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[20]^u[18]^u[17]^u[15]^u[13]^u[11]^u[8]^u[7]^u[6]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[280] = x[248]^x[298]^x[299]^x[300]^x[303]^x[305]^x[312]^x[313]^x[315]^x[316]^x[317]^x[318]^x[320]^x[322]^x[327]^x[328]^x[329]^u[31]^u[30]^u[29]^u[26]^u[24]^u[17]^u[16]^u[14]^u[13]^u[12]^u[11]^u[9]^u[7]^u[2]^u[1]^u[0];
	y[281] = x[249]^x[298]^x[302]^x[307]^x[310]^x[313]^x[314]^x[317]^x[320]^x[321]^x[324]^x[325]^x[326]^x[327]^x[328]^x[329]^u[31]^u[27]^u[22]^u[19]^u[16]^u[15]^u[12]^u[9]^u[8]^u[5]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[282] = x[250]^x[298]^x[300]^x[301]^x[302]^x[303]^x[304]^x[306]^x[307]^x[308]^x[310]^x[311]^x[314]^x[315]^x[316]^x[319]^x[320]^x[321]^x[322]^x[323]^x[324]^x[328]^x[329]^u[31]^u[29]^u[28]^u[27]^u[26]^u[25]^u[23]^u[22]^u[21]^u[19]^u[18]^u[15]^u[14]^u[13]^u[10]^u[9]^u[8]^u[7]^u[6]^u[5]^u[1]^u[0];
	y[283] = x[251]^x[299]^x[301]^x[302]^x[303]^x[304]^x[305]^x[307]^x[308]^x[309]^x[311]^x[312]^x[315]^x[316]^x[317]^x[320]^x[321]^x[322]^x[323]^x[324]^x[325]^x[329]^u[30]^u[28]^u[27]^u[26]^u[25]^u[24]^u[22]^u[21]^u[20]^u[18]^u[17]^u[14]^u[13]^u[12]^u[9]^u[8]^u[7]^u[6]^u[5]^u[4]^u[0];
	y[284] = x[252]^x[298]^x[299]^x[301]^x[303]^x[305]^x[307]^x[308]^x[309]^x[312]^x[313]^x[317]^x[319]^x[320]^x[321]^x[322]^x[327]^u[31]^u[30]^u[28]^u[26]^u[24]^u[22]^u[21]^u[20]^u[17]^u[16]^u[12]^u[10]^u[9]^u[8]^u[7]^u[2];
	y[285] = x[253]^x[298]^x[301]^x[307]^x[308]^x[309]^x[313]^x[314]^x[316]^x[319]^x[321]^x[322]^x[324]^x[325]^x[326]^x[327]^x[328]^u[31]^u[28]^u[22]^u[21]^u[20]^u[16]^u[15]^u[13]^u[10]^u[8]^u[7]^u[5]^u[4]^u[3]^u[2]^u[1];
	y[286] = x[254]^x[299]^x[302]^x[308]^x[309]^x[310]^x[314]^x[315]^x[317]^x[320]^x[322]^x[323]^x[325]^x[326]^x[327]^x[328]^x[329]^u[30]^u[27]^u[21]^u[20]^u[19]^u[15]^u[14]^u[12]^u[9]^u[7]^u[6]^u[4]^u[3]^u[2]^u[1]^u[0];
	y[287] = x[255]^x[298]^x[299]^x[301]^x[302]^x[303]^x[304]^x[306]^x[307]^x[309]^x[311]^x[315]^x[319]^x[320]^x[321]^x[325]^x[328]^x[329]^u[31]^u[30]^u[28]^u[27]^u[26]^u[25]^u[23]^u[22]^u[20]^u[18]^u[14]^u[10]^u[9]^u[8]^u[4]^u[1]^u[0];
	y[288] = x[256]^x[299]^x[300]^x[302]^x[303]^x[304]^x[305]^x[307]^x[308]^x[310]^x[312]^x[316]^x[320]^x[321]^x[322]^x[326]^x[329]^u[30]^u[29]^u[27]^u[26]^u[25]^u[24]^u[22]^u[21]^u[19]^u[17]^u[13]^u[9]^u[8]^u[7]^u[3]^u[0];
	y[289] = x[257]^x[298]^x[299]^x[302]^x[303]^x[305]^x[307]^x[308]^x[309]^x[310]^x[311]^x[313]^x[316]^x[317]^x[318]^x[319]^x[320]^x[321]^x[322]^x[324]^x[325]^x[326]^u[31]^u[30]^u[27]^u[26]^u[24]^u[22]^u[21]^u[20]^u[19]^u[18]^u[16]^u[13]^u[12]^u[11]^u[10]^u[9]^u[8]^u[7]^u[5]^u[4]^u[3];
	y[290] = x[258]^x[298]^x[301]^x[302]^x[303]^x[307]^x[308]^x[309]^x[311]^x[312]^x[314]^x[316]^x[317]^x[321]^x[322]^x[324]^u[31]^u[28]^u[27]^u[26]^u[22]^u[21]^u[20]^u[18]^u[17]^u[15]^u[13]^u[12]^u[8]^u[7]^u[5];
	y[291] = x[259]^x[299]^x[302]^x[303]^x[304]^x[308]^x[309]^x[310]^x[312]^x[313]^x[315]^x[317]^x[318]^x[322]^x[323]^x[325]^u[30]^u[27]^u[26]^u[25]^u[21]^u[20]^u[19]^u[17]^u[16]^u[14]^u[12]^u[11]^u[7]^u[6]^u[4];
	y[292] = x[260]^x[300]^x[303]^x[304]^x[305]^x[309]^x[310]^x[311]^x[313]^x[314]^x[316]^x[318]^x[319]^x[323]^x[324]^x[326]^u[29]^u[26]^u[25]^u[24]^u[20]^u[19]^u[18]^u[16]^u[15]^u[13]^u[11]^u[10]^u[6]^u[5]^u[3];
	y[293] = x[261]^x[298]^x[299]^x[300]^x[302]^x[305]^x[307]^x[311]^x[312]^x[314]^x[315]^x[316]^x[317]^x[318]^x[323]^x[326]^u[31]^u[30]^u[29]^u[27]^u[24]^u[22]^u[18]^u[17]^u[15]^u[14]^u[13]^u[12]^u[11]^u[6]^u[3];
	y[294] = x[262]^x[299]^x[300]^x[301]^x[303]^x[306]^x[308]^x[312]^x[313]^x[315]^x[316]^x[317]^x[318]^x[319]^x[324]^x[327]^u[30]^u[29]^u[28]^u[26]^u[23]^u[21]^u[17]^u[16]^u[14]^u[13]^u[12]^u[11]^u[10]^u[5]^u[2];
	y[295] = x[263]^x[298]^x[299]^x[306]^x[309]^x[310]^x[313]^x[314]^x[317]^x[323]^x[324]^x[326]^x[327]^x[328]^u[31]^u[30]^u[23]^u[20]^u[19]^u[16]^u[15]^u[12]^u[6]^u[5]^u[3]^u[2]^u[1];
	y[296] = x[264]^x[299]^x[300]^x[307]^x[310]^x[311]^x[314]^x[315]^x[318]^x[324]^x[325]^x[327]^x[328]^x[329]^u[30]^u[29]^u[22]^u[19]^u[18]^u[15]^u[14]^u[11]^u[5]^u[4]^u[2]^u[1]^u[0];
	y[297] = x[265]^x[298]^x[299]^x[302]^x[304]^x[306]^x[307]^x[308]^x[310]^x[311]^x[312]^x[315]^x[318]^x[320]^x[323]^x[324]^x[327]^x[328]^x[329]^u[31]^u[30]^u[27]^u[25]^u[23]^u[22]^u[21]^u[19]^u[18]^u[17]^u[14]^u[11]^u[9]^u[6]^u[5]^u[2]^u[1]^u[0];
	y[298] = x[266]^x[298]^x[301]^x[302]^x[303]^x[304]^x[305]^x[306]^x[308]^x[309]^x[310]^x[311]^x[312]^x[313]^x[318]^x[320]^x[321]^x[323]^x[326]^x[327]^x[328]^x[329]^u[31]^u[28]^u[27]^u[26]^u[25]^u[24]^u[23]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[11]^u[9]^u[8]^u[6]^u[3]^u[2]^u[1]^u[0];
	y[299] = x[267]^x[299]^x[302]^x[303]^x[304]^x[305]^x[306]^x[307]^x[309]^x[310]^x[311]^x[312]^x[313]^x[314]^x[319]^x[321]^x[322]^x[324]^x[327]^x[328]^x[329]^u[30]^u[27]^u[26]^u[25]^u[24]^u[23]^u[22]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[10]^u[8]^u[7]^u[5]^u[2]^u[1]^u[0];
	y[300] = x[268]^x[300]^x[303]^x[304]^x[305]^x[306]^x[307]^x[308]^x[310]^x[311]^x[312]^x[313]^x[314]^x[315]^x[320]^x[322]^x[323]^x[325]^x[328]^x[329]^u[29]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[9]^u[7]^u[6]^u[4]^u[1]^u[0];
	y[301] = x[269]^x[298]^x[299]^x[300]^x[302]^x[305]^x[308]^x[309]^x[310]^x[311]^x[312]^x[313]^x[314]^x[315]^x[318]^x[319]^x[320]^x[321]^x[325]^x[327]^x[329]^u[31]^u[30]^u[29]^u[27]^u[24]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[11]^u[10]^u[9]^u[8]^u[4]^u[2]^u[0];
	y[302] = x[270]^x[299]^x[300]^x[301]^x[303]^x[306]^x[309]^x[310]^x[311]^x[312]^x[313]^x[314]^x[315]^x[316]^x[319]^x[320]^x[321]^x[322]^x[326]^x[328]^u[30]^u[29]^u[28]^u[26]^u[23]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[13]^u[10]^u[9]^u[8]^u[7]^u[3]^u[1];
	y[303] = x[271]^x[300]^x[301]^x[302]^x[304]^x[307]^x[310]^x[311]^x[312]^x[313]^x[314]^x[315]^x[316]^x[317]^x[320]^x[321]^x[322]^x[323]^x[327]^x[329]^u[29]^u[28]^u[27]^u[25]^u[22]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[13]^u[12]^u[9]^u[8]^u[7]^u[6]^u[2]^u[0];
	y[304] = x[272]^x[298]^x[299]^x[300]^x[303]^x[304]^x[305]^x[306]^x[307]^x[308]^x[310]^x[311]^x[312]^x[313]^x[314]^x[315]^x[317]^x[319]^x[320]^x[321]^x[322]^x[325]^x[326]^x[327]^x[328]^u[31]^u[30]^u[29]^u[26]^u[25]^u[24]^u[23]^u[22]^u[21]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[10]^u[9]^u[8]^u[7]^u[4]^u[3]^u[2]^u[1];
	y[305] = x[273]^x[298]^x[302]^x[305]^x[308]^x[309]^x[310]^x[311]^x[312]^x[313]^x[314]^x[315]^x[319]^x[321]^x[322]^x[324]^x[325]^x[328]^x[329]^u[31]^u[27]^u[24]^u[21]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[10]^u[8]^u[7]^u[5]^u[4]^u[1]^u[0];
	y[306] = x[274]^x[299]^x[303]^x[306]^x[309]^x[310]^x[311]^x[312]^x[313]^x[314]^x[315]^x[316]^x[320]^x[322]^x[323]^x[325]^x[326]^x[329]^u[30]^u[26]^u[23]^u[20]^u[19]^u[18]^u[17]^u[16]^u[15]^u[14]^u[13]^u[9]^u[7]^u[6]^u[4]^u[3]^u[0];
	y[307] = x[275]^x[298]^x[299]^x[301]^x[302]^x[306]^x[311]^x[312]^x[313]^x[314]^x[315]^x[317]^x[318]^x[319]^x[320]^x[321]^x[325]^u[31]^u[30]^u[28]^u[27]^u[23]^u[18]^u[17]^u[16]^u[15]^u[14]^u[12]^u[11]^u[10]^u[9]^u[8]^u[4];
	y[308] = x[276]^x[299]^x[300]^x[302]^x[303]^x[307]^x[312]^x[313]^x[314]^x[315]^x[316]^x[318]^x[319]^x[320]^x[321]^x[322]^x[326]^u[30]^u[29]^u[27]^u[26]^u[22]^u[17]^u[16]^u[15]^u[14]^u[13]^u[11]^u[10]^u[9]^u[8]^u[7]^u[3];
	y[309] = x[277]^x[300]^x[301]^x[303]^x[304]^x[308]^x[313]^x[314]^x[315]^x[316]^x[317]^x[319]^x[320]^x[321]^x[322]^x[323]^x[327]^u[29]^u[28]^u[26]^u[25]^u[21]^u[16]^u[15]^u[14]^u[13]^u[12]^u[10]^u[9]^u[8]^u[7]^u[6]^u[2];
	y[310] = x[278]^x[298]^x[299]^x[300]^x[305]^x[306]^x[307]^x[309]^x[310]^x[314]^x[315]^x[317]^x[319]^x[321]^x[322]^x[325]^x[326]^x[327]^x[328]^u[31]^u[30]^u[29]^u[24]^u[23]^u[22]^u[20]^u[19]^u[15]^u[14]^u[12]^u[10]^u[8]^u[7]^u[4]^u[3]^u[2]^u[1];
	y[311] = x[279]^x[299]^x[300]^x[301]^x[306]^x[307]^x[308]^x[310]^x[311]^x[315]^x[316]^x[318]^x[320]^x[322]^x[323]^x[326]^x[327]^x[328]^x[329]^u[30]^u[29]^u[28]^u[23]^u[22]^u[21]^u[19]^u[18]^u[14]^u[13]^u[11]^u[9]^u[7]^u[6]^u[3]^u[2]^u[1]^u[0];
	y[312] = x[280]^x[298]^x[299]^x[304]^x[306]^x[308]^x[309]^x[310]^x[311]^x[312]^x[317]^x[318]^x[320]^x[321]^x[325]^x[326]^x[328]^x[329]^u[31]^u[30]^u[25]^u[23]^u[21]^u[20]^u[19]^u[18]^u[17]^u[12]^u[11]^u[9]^u[8]^u[4]^u[3]^u[1]^u[0];
	y[313] = x[281]^x[299]^x[300]^x[305]^x[307]^x[309]^x[310]^x[311]^x[312]^x[313]^x[318]^x[319]^x[321]^x[322]^x[326]^x[327]^x[329]^u[30]^u[29]^u[24]^u[22]^u[20]^u[19]^u[18]^u[17]^u[16]^u[11]^u[10]^u[8]^u[7]^u[3]^u[2]^u[0];
	y[314] = x[282]^x[298]^x[299]^x[302]^x[304]^x[307]^x[308]^x[311]^x[312]^x[313]^x[314]^x[316]^x[318]^x[322]^x[324]^x[325]^x[326]^x[328]^u[31]^u[30]^u[27]^u[25]^u[22]^u[21]^u[18]^u[17]^u[16]^u[15]^u[13]^u[11]^u[7]^u[5]^u[4]^u[3]^u[1];
	y[315] = x[283]^x[299]^x[300]^x[303]^x[305]^x[308]^x[309]^x[312]^x[313]^x[314]^x[315]^x[317]^x[319]^x[323]^x[325]^x[326]^x[327]^x[329]^u[30]^u[29]^u[26]^u[24]^u[21]^u[20]^u[17]^u[16]^u[15]^u[14]^u[12]^u[10]^u[6]^u[4]^u[3]^u[2]^u[0];
	y[316] = x[284]^x[300]^x[301]^x[304]^x[306]^x[309]^x[310]^x[313]^x[314]^x[315]^x[316]^x[318]^x[320]^x[324]^x[326]^x[327]^x[328]^u[29]^u[28]^u[25]^u[23]^u[20]^u[19]^u[16]^u[15]^u[14]^u[13]^u[11]^u[9]^u[5]^u[3]^u[2]^u[1];
	y[317] = x[285]^x[298]^x[299]^x[300]^x[304]^x[305]^x[306]^x[311]^x[314]^x[315]^x[317]^x[318]^x[320]^x[321]^x[323]^x[324]^x[326]^x[328]^x[329]^u[31]^u[30]^u[29]^u[25]^u[24]^u[23]^u[18]^u[15]^u[14]^u[12]^u[11]^u[9]^u[8]^u[6]^u[5]^u[3]^u[1]^u[0];
	y[318] = x[286]^x[299]^x[300]^x[301]^x[305]^x[306]^x[307]^x[312]^x[315]^x[316]^x[318]^x[319]^x[321]^x[322]^x[324]^x[325]^x[327]^x[329]^u[30]^u[29]^u[28]^u[24]^u[23]^u[22]^u[17]^u[14]^u[13]^u[11]^u[10]^u[8]^u[7]^u[5]^u[4]^u[2]^u[0];
	y[319] = x[287]^x[300]^x[301]^x[302]^x[306]^x[307]^x[308]^x[313]^x[316]^x[317]^x[319]^x[320]^x[322]^x[323]^x[325]^x[326]^x[328]^u[29]^u[28]^u[27]^u[23]^u[22]^u[21]^u[16]^u[13]^u[12]^u[10]^u[9]^u[7]^u[6]^u[4]^u[3]^u[1];
	y[320] = x[288]^x[301]^x[302]^x[303]^x[307]^x[308]^x[309]^x[314]^x[317]^x[318]^x[320]^x[321]^x[323]^x[324]^x[326]^x[327]^x[329]^u[28]^u[27]^u[26]^u[22]^u[21]^u[20]^u[15]^u[12]^u[11]^u[9]^u[8]^u[6]^u[5]^u[3]^u[2]^u[0];
	y[321] = x[289]^x[298]^x[299]^x[300]^x[301]^x[303]^x[306]^x[307]^x[308]^x[309]^x[315]^x[316]^x[320]^x[321]^x[322]^x[323]^x[326]^x[328]^u[31]^u[30]^u[29]^u[28]^u[26]^u[23]^u[22]^u[21]^u[20]^u[14]^u[13]^u[9]^u[8]^u[7]^u[6]^u[3]^u[1];
	y[322] = x[290]^x[299]^x[300]^x[301]^x[302]^x[304]^x[307]^x[308]^x[309]^x[310]^x[316]^x[317]^x[321]^x[322]^x[323]^x[324]^x[327]^x[329]^u[30]^u[29]^u[28]^u[27]^u[25]^u[22]^u[21]^u[20]^u[19]^u[13]^u[12]^u[8]^u[7]^u[6]^u[5]^u[2]^u[0];
	y[323] = x[291]^x[300]^x[301]^x[302]^x[303]^x[305]^x[308]^x[309]^x[310]^x[311]^x[317]^x[318]^x[322]^x[323]^x[324]^x[325]^x[328]^u[29]^u[28]^u[27]^u[26]^u[24]^u[21]^u[20]^u[19]^u[18]^u[12]^u[11]^u[7]^u[6]^u[5]^u[4]^u[1];
	y[324] = x[292]^x[301]^x[302]^x[303]^x[304]^x[306]^x[309]^x[310]^x[311]^x[312]^x[318]^x[319]^x[323]^x[324]^x[325]^x[326]^x[329]^u[28]^u[27]^u[26]^u[25]^u[23]^u[20]^u[19]^u[18]^u[17]^u[11]^u[10]^u[6]^u[5]^u[4]^u[3]^u[0];
	y[325] = x[293]^x[298]^x[299]^x[300]^x[301]^x[303]^x[305]^x[306]^x[311]^x[312]^x[313]^x[316]^x[318]^x[323]^u[31]^u[30]^u[29]^u[28]^u[26]^u[24]^u[23]^u[18]^u[17]^u[16]^u[13]^u[11]^u[6];
	y[326] = x[294]^x[299]^x[300]^x[301]^x[302]^x[304]^x[306]^x[307]^x[312]^x[313]^x[314]^x[317]^x[319]^x[324]^u[30]^u[29]^u[28]^u[27]^u[25]^u[23]^u[22]^u[17]^u[16]^u[15]^u[12]^u[10]^u[5];
	y[327] = x[295]^x[300]^x[301]^x[302]^x[303]^x[305]^x[307]^x[308]^x[313]^x[314]^x[315]^x[318]^x[320]^x[325]^u[29]^u[28]^u[27]^u[26]^u[24]^u[22]^u[21]^u[16]^u[15]^u[14]^u[11]^u[9]^u[4];
	y[328] = x[296]^x[301]^x[302]^x[303]^x[304]^x[306]^x[308]^x[309]^x[314]^x[315]^x[316]^x[319]^x[321]^x[326]^u[28]^u[27]^u[26]^u[25]^u[23]^u[21]^u[20]^u[15]^u[14]^u[13]^u[10]^u[8]^u[3];
	y[329] = x[297]^x[298]^x[299]^x[300]^x[301]^x[303]^x[305]^x[306]^x[309]^x[315]^x[317]^x[318]^x[319]^x[322]^x[323]^x[324]^x[325]^x[326]^u[31]^u[30]^u[29]^u[28]^u[26]^u[24]^u[23]^u[20]^u[14]^u[12]^u[11]^u[10]^u[7]^u[6]^u[5]^u[4]^u[3];
	return y;
endfunction
