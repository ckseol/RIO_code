package RS_common;
import Vector::*;

typedef Bit#(6) SYMBOL;
typedef 63 CODEWORD_LEN;
typedef Vector#(18, SYMBOL) SYNDROME;
typedef 6 SYM_CNT_BIT_WIDTH;

typedef 9 T_RS;
typedef 18 DOUBLE_T_RS;
typedef Vector#(19, SYMBOL) POLYNOMIAL;
typedef UInt#(8) POLY_IDX;

typedef 45 MESSAGE_LEN;
typedef 18  PARITY_LEN;
typedef Vector#(18, SYMBOL) PARITY;


(* noinline *)
function Bit#(6) gf_mul_m6(Bit#(6) a, Bit#(6) b);
        Bit#(6) c;
        Bit#(11) c_tmp;
        c_tmp[0] = (a[0] & b[0]);
        c_tmp[1] = (a[0] & b[1])^(a[1] & b[0]);
        c_tmp[2] = (a[0] & b[2])^(a[1] & b[1])^(a[2] & b[0]);
        c_tmp[3] = (a[0] & b[3])^(a[1] & b[2])^(a[2] & b[1])^(a[3] & b[0]);
        c_tmp[4] = (a[0] & b[4])^(a[1] & b[3])^(a[2] & b[2])^(a[3] & b[1])^(a[4] & b[0]);
        c_tmp[5] = (a[0] & b[5])^(a[1] & b[4])^(a[2] & b[3])^(a[3] & b[2])^(a[4] & b[1])^(a[5] & b[0]);
        c_tmp[6] = (a[1] & b[5])^(a[2] & b[4])^(a[3] & b[3])^(a[4] & b[2])^(a[5] & b[1]);
        c_tmp[7] = (a[2] & b[5])^(a[3] & b[4])^(a[4] & b[3])^(a[5] & b[2]);
        c_tmp[8] = (a[3] & b[5])^(a[4] & b[4])^(a[5] & b[3]);
        c_tmp[9] = (a[4] & b[5])^(a[5] & b[4]);
        c_tmp[10] = (a[5] & b[5]);
        c[0] = c_tmp[0]^c_tmp[6];
        c[1] = c_tmp[1]^c_tmp[6]^c_tmp[7];
        c[2] = c_tmp[2]^c_tmp[7]^c_tmp[8];
        c[3] = c_tmp[3]^c_tmp[8]^c_tmp[9];
        c[4] = c_tmp[4]^c_tmp[9]^c_tmp[10];
        c[5] = c_tmp[5]^c_tmp[10];
        return c;
endfunction

(* noinline *)
function Vector#(18, Bit#(6)) get_alpha_list(UInt#(6) loc_j);
	Vector#(18, Bit#(6)) a = replicate(0);
	case(loc_j)
	6'd0 : begin a[0]=6'd1; a[1]=6'd1; a[2]=6'd1; a[3]=6'd1; a[4]=6'd1; a[5]=6'd1; a[6]=6'd1; a[7]=6'd1; a[8]=6'd1; a[9]=6'd1; a[10]=6'd1; a[11]=6'd1; a[12]=6'd1; a[13]=6'd1; a[14]=6'd1; a[15]=6'd1; a[16]=6'd1; a[17]=6'd1;  end
	6'd1 : begin a[0]=6'd33; a[1]=6'd49; a[2]=6'd57; a[3]=6'd61; a[4]=6'd63; a[5]=6'd62; a[6]=6'd31; a[7]=6'd46; a[8]=6'd23; a[9]=6'd42; a[10]=6'd21; a[11]=6'd43; a[12]=6'd52; a[13]=6'd26; a[14]=6'd13; a[15]=6'd39; a[16]=6'd50; a[17]=6'd25;  end
	6'd2 : begin a[0]=6'd49; a[1]=6'd61; a[2]=6'd62; a[3]=6'd46; a[4]=6'd42; a[5]=6'd43; a[6]=6'd26; a[7]=6'd39; a[8]=6'd25; a[9]=6'd55; a[10]=6'd29; a[11]=6'd54; a[12]=6'd44; a[13]=6'd11; a[14]=6'd18; a[15]=6'd37; a[16]=6'd56; a[17]=6'd14;  end
	6'd3 : begin a[0]=6'd57; a[1]=6'd62; a[2]=6'd23; a[3]=6'd43; a[4]=6'd13; a[5]=6'd25; a[6]=6'd58; a[7]=6'd54; a[8]=6'd22; a[9]=6'd18; a[10]=6'd51; a[11]=6'd14; a[12]=6'd17; a[13]=6'd59; a[14]=6'd15; a[15]=6'd40; a[16]=6'd5; a[17]=6'd24;  end
	6'd4 : begin a[0]=6'd61; a[1]=6'd46; a[2]=6'd43; a[3]=6'd39; a[4]=6'd55; a[5]=6'd54; a[6]=6'd11; a[7]=6'd37; a[8]=6'd14; a[9]=6'd41; a[10]=6'd30; a[11]=6'd40; a[12]=6'd35; a[13]=6'd6; a[14]=6'd8; a[15]=6'd33; a[16]=6'd63; a[17]=6'd23;  end
	6'd5 : begin a[0]=6'd63; a[1]=6'd42; a[2]=6'd13; a[3]=6'd55; a[4]=6'd27; a[5]=6'd18; a[6]=6'd28; a[7]=6'd41; a[8]=6'd15; a[9]=6'd10; a[10]=6'd12; a[11]=6'd8; a[12]=6'd49; a[13]=6'd31; a[14]=6'd43; a[15]=6'd50; a[16]=6'd29; a[17]=6'd22;  end
	6'd6 : begin a[0]=6'd62; a[1]=6'd43; a[2]=6'd25; a[3]=6'd54; a[4]=6'd18; a[5]=6'd14; a[6]=6'd59; a[7]=6'd40; a[8]=6'd24; a[9]=6'd8; a[10]=6'd57; a[11]=6'd23; a[12]=6'd13; a[13]=6'd58; a[14]=6'd22; a[15]=6'd51; a[16]=6'd17; a[17]=6'd15;  end
	6'd7 : begin a[0]=6'd31; a[1]=6'd26; a[2]=6'd58; a[3]=6'd11; a[4]=6'd28; a[5]=6'd59; a[6]=6'd20; a[7]=6'd6; a[8]=6'd1; a[9]=6'd31; a[10]=6'd26; a[11]=6'd58; a[12]=6'd11; a[13]=6'd28; a[14]=6'd59; a[15]=6'd20; a[16]=6'd6; a[17]=6'd1;  end
	6'd8 : begin a[0]=6'd46; a[1]=6'd39; a[2]=6'd54; a[3]=6'd37; a[4]=6'd41; a[5]=6'd40; a[6]=6'd6; a[7]=6'd33; a[8]=6'd23; a[9]=6'd50; a[10]=6'd27; a[11]=6'd51; a[12]=6'd53; a[13]=6'd20; a[14]=6'd3; a[15]=6'd49; a[16]=6'd42; a[17]=6'd25;  end
	6'd9 : begin a[0]=6'd23; a[1]=6'd25; a[2]=6'd22; a[3]=6'd14; a[4]=6'd15; a[5]=6'd24; a[6]=6'd1; a[7]=6'd23; a[8]=6'd25; a[9]=6'd22; a[10]=6'd14; a[11]=6'd15; a[12]=6'd24; a[13]=6'd1; a[14]=6'd23; a[15]=6'd25; a[16]=6'd22; a[17]=6'd14;  end
	6'd10 : begin a[0]=6'd42; a[1]=6'd55; a[2]=6'd18; a[3]=6'd41; a[4]=6'd10; a[5]=6'd8; a[6]=6'd31; a[7]=6'd50; a[8]=6'd22; a[9]=6'd7; a[10]=6'd19; a[11]=6'd3; a[12]=6'd61; a[13]=6'd26; a[14]=6'd54; a[15]=6'd56; a[16]=6'd30; a[17]=6'd24;  end
	6'd11 : begin a[0]=6'd21; a[1]=6'd29; a[2]=6'd51; a[3]=6'd30; a[4]=6'd12; a[5]=6'd57; a[6]=6'd26; a[7]=6'd27; a[8]=6'd14; a[9]=6'd19; a[10]=6'd32; a[11]=6'd62; a[12]=6'd50; a[13]=6'd11; a[14]=6'd17; a[15]=6'd10; a[16]=6'd4; a[17]=6'd23;  end
	6'd12 : begin a[0]=6'd43; a[1]=6'd54; a[2]=6'd14; a[3]=6'd40; a[4]=6'd8; a[5]=6'd23; a[6]=6'd58; a[7]=6'd51; a[8]=6'd15; a[9]=6'd3; a[10]=6'd62; a[11]=6'd25; a[12]=6'd18; a[13]=6'd59; a[14]=6'd24; a[15]=6'd57; a[16]=6'd13; a[17]=6'd22;  end
	6'd13 : begin a[0]=6'd52; a[1]=6'd44; a[2]=6'd17; a[3]=6'd35; a[4]=6'd49; a[5]=6'd13; a[6]=6'd11; a[7]=6'd53; a[8]=6'd24; a[9]=6'd61; a[10]=6'd50; a[11]=6'd18; a[12]=6'd60; a[13]=6'd6; a[14]=6'd62; a[15]=6'd45; a[16]=6'd37; a[17]=6'd15;  end
	6'd14 : begin a[0]=6'd26; a[1]=6'd11; a[2]=6'd59; a[3]=6'd6; a[4]=6'd31; a[5]=6'd58; a[6]=6'd28; a[7]=6'd20; a[8]=6'd1; a[9]=6'd26; a[10]=6'd11; a[11]=6'd59; a[12]=6'd6; a[13]=6'd31; a[14]=6'd58; a[15]=6'd28; a[16]=6'd20; a[17]=6'd1;  end
	6'd15 : begin a[0]=6'd13; a[1]=6'd18; a[2]=6'd15; a[3]=6'd8; a[4]=6'd43; a[5]=6'd22; a[6]=6'd59; a[7]=6'd3; a[8]=6'd23; a[9]=6'd54; a[10]=6'd17; a[11]=6'd24; a[12]=6'd62; a[13]=6'd58; a[14]=6'd14; a[15]=6'd5; a[16]=6'd57; a[17]=6'd25;  end
	6'd16 : begin a[0]=6'd39; a[1]=6'd37; a[2]=6'd40; a[3]=6'd33; a[4]=6'd50; a[5]=6'd51; a[6]=6'd20; a[7]=6'd49; a[8]=6'd25; a[9]=6'd56; a[10]=6'd10; a[11]=6'd57; a[12]=6'd45; a[13]=6'd28; a[14]=6'd5; a[15]=6'd61; a[16]=6'd55; a[17]=6'd14;  end
	6'd17 : begin a[0]=6'd50; a[1]=6'd56; a[2]=6'd5; a[3]=6'd63; a[4]=6'd29; a[5]=6'd17; a[6]=6'd6; a[7]=6'd42; a[8]=6'd22; a[9]=6'd30; a[10]=6'd4; a[11]=6'd13; a[12]=6'd37; a[13]=6'd20; a[14]=6'd57; a[15]=6'd55; a[16]=6'd7; a[17]=6'd24;  end
	6'd18 : begin a[0]=6'd25; a[1]=6'd14; a[2]=6'd24; a[3]=6'd23; a[4]=6'd22; a[5]=6'd15; a[6]=6'd1; a[7]=6'd25; a[8]=6'd14; a[9]=6'd24; a[10]=6'd23; a[11]=6'd22; a[12]=6'd15; a[13]=6'd1; a[14]=6'd25; a[15]=6'd14; a[16]=6'd24; a[17]=6'd23;  end
	6'd19 : begin a[0]=6'd45; a[1]=6'd34; a[2]=6'd3; a[3]=6'd52; a[4]=6'd37; a[5]=6'd5; a[6]=6'd31; a[7]=6'd44; a[8]=6'd15; a[9]=6'd33; a[10]=6'd55; a[11]=6'd17; a[12]=6'd32; a[13]=6'd26; a[14]=6'd51; a[15]=6'd35; a[16]=6'd46; a[17]=6'd22;  end
	6'd20 : begin a[0]=6'd55; a[1]=6'd41; a[2]=6'd8; a[3]=6'd50; a[4]=6'd7; a[5]=6'd3; a[6]=6'd26; a[7]=6'd56; a[8]=6'd24; a[9]=6'd21; a[10]=6'd9; a[11]=6'd5; a[12]=6'd46; a[13]=6'd11; a[14]=6'd40; a[15]=6'd63; a[16]=6'd27; a[17]=6'd15;  end
	6'd21 : begin a[0]=6'd58; a[1]=6'd59; a[2]=6'd1; a[3]=6'd58; a[4]=6'd59; a[5]=6'd1; a[6]=6'd58; a[7]=6'd59; a[8]=6'd1; a[9]=6'd58; a[10]=6'd59; a[11]=6'd1; a[12]=6'd58; a[13]=6'd59; a[14]=6'd1; a[15]=6'd58; a[16]=6'd59; a[17]=6'd1;  end
	6'd22 : begin a[0]=6'd29; a[1]=6'd30; a[2]=6'd57; a[3]=6'd27; a[4]=6'd19; a[5]=6'd62; a[6]=6'd11; a[7]=6'd10; a[8]=6'd23; a[9]=6'd9; a[10]=6'd48; a[11]=6'd43; a[12]=6'd56; a[13]=6'd6; a[14]=6'd13; a[15]=6'd7; a[16]=6'd16; a[17]=6'd25;  end
	6'd23 : begin a[0]=6'd47; a[1]=6'd38; a[2]=6'd62; a[3]=6'd36; a[4]=6'd35; a[5]=6'd43; a[6]=6'd28; a[7]=6'd32; a[8]=6'd25; a[9]=6'd53; a[10]=6'd33; a[11]=6'd54; a[12]=6'd19; a[13]=6'd31; a[14]=6'd18; a[15]=6'd48; a[16]=6'd52; a[17]=6'd14;  end
	6'd24 : begin a[0]=6'd54; a[1]=6'd40; a[2]=6'd23; a[3]=6'd51; a[4]=6'd3; a[5]=6'd25; a[6]=6'd59; a[7]=6'd57; a[8]=6'd22; a[9]=6'd5; a[10]=6'd43; a[11]=6'd14; a[12]=6'd8; a[13]=6'd58; a[14]=6'd15; a[15]=6'd62; a[16]=6'd18; a[17]=6'd24;  end
	6'd25 : begin a[0]=6'd27; a[1]=6'd10; a[2]=6'd43; a[3]=6'd7; a[4]=6'd2; a[5]=6'd54; a[6]=6'd20; a[7]=6'd21; a[8]=6'd14; a[9]=6'd4; a[10]=6'd47; a[11]=6'd40; a[12]=6'd42; a[13]=6'd28; a[14]=6'd8; a[15]=6'd29; a[16]=6'd19; a[17]=6'd23;  end
	6'd26 : begin a[0]=6'd44; a[1]=6'd35; a[2]=6'd13; a[3]=6'd53; a[4]=6'd61; a[5]=6'd18; a[6]=6'd6; a[7]=6'd45; a[8]=6'd15; a[9]=6'd46; a[10]=6'd56; a[11]=6'd8; a[12]=6'd47; a[13]=6'd20; a[14]=6'd43; a[15]=6'd34; a[16]=6'd33; a[17]=6'd22;  end
	6'd27 : begin a[0]=6'd22; a[1]=6'd24; a[2]=6'd25; a[3]=6'd15; a[4]=6'd23; a[5]=6'd14; a[6]=6'd1; a[7]=6'd22; a[8]=6'd24; a[9]=6'd25; a[10]=6'd15; a[11]=6'd23; a[12]=6'd14; a[13]=6'd1; a[14]=6'd22; a[15]=6'd24; a[16]=6'd25; a[17]=6'd15;  end
	6'd28 : begin a[0]=6'd11; a[1]=6'd6; a[2]=6'd58; a[3]=6'd20; a[4]=6'd26; a[5]=6'd59; a[6]=6'd31; a[7]=6'd28; a[8]=6'd1; a[9]=6'd11; a[10]=6'd6; a[11]=6'd58; a[12]=6'd20; a[13]=6'd26; a[14]=6'd59; a[15]=6'd31; a[16]=6'd28; a[17]=6'd1;  end
	6'd29 : begin a[0]=6'd36; a[1]=6'd32; a[2]=6'd54; a[3]=6'd48; a[4]=6'd45; a[5]=6'd40; a[6]=6'd26; a[7]=6'd60; a[8]=6'd23; a[9]=6'd34; a[10]=6'd61; a[11]=6'd51; a[12]=6'd2; a[13]=6'd11; a[14]=6'd3; a[15]=6'd47; a[16]=6'd35; a[17]=6'd25;  end
	6'd30 : begin a[0]=6'd18; a[1]=6'd8; a[2]=6'd22; a[3]=6'd3; a[4]=6'd54; a[5]=6'd24; a[6]=6'd58; a[7]=6'd5; a[8]=6'd25; a[9]=6'd40; a[10]=6'd13; a[11]=6'd15; a[12]=6'd43; a[13]=6'd59; a[14]=6'd23; a[15]=6'd17; a[16]=6'd62; a[17]=6'd14;  end
	6'd31 : begin a[0]=6'd9; a[1]=6'd2; a[2]=6'd18; a[3]=6'd4; a[4]=6'd36; a[5]=6'd8; a[6]=6'd11; a[7]=6'd16; a[8]=6'd22; a[9]=6'd32; a[10]=6'd44; a[11]=6'd3; a[12]=6'd27; a[13]=6'd6; a[14]=6'd54; a[15]=6'd12; a[16]=6'd47; a[17]=6'd24;  end
	6'd32 : begin a[0]=6'd37; a[1]=6'd33; a[2]=6'd51; a[3]=6'd49; a[4]=6'd56; a[5]=6'd57; a[6]=6'd28; a[7]=6'd61; a[8]=6'd14; a[9]=6'd63; a[10]=6'd7; a[11]=6'd62; a[12]=6'd34; a[13]=6'd31; a[14]=6'd17; a[15]=6'd46; a[16]=6'd41; a[17]=6'd23;  end
	6'd33 : begin a[0]=6'd51; a[1]=6'd57; a[2]=6'd14; a[3]=6'd62; a[4]=6'd17; a[5]=6'd23; a[6]=6'd59; a[7]=6'd43; a[8]=6'd15; a[9]=6'd13; a[10]=6'd40; a[11]=6'd25; a[12]=6'd5; a[13]=6'd58; a[14]=6'd24; a[15]=6'd54; a[16]=6'd3; a[17]=6'd22;  end
	6'd34 : begin a[0]=6'd56; a[1]=6'd63; a[2]=6'd17; a[3]=6'd42; a[4]=6'd30; a[5]=6'd13; a[6]=6'd20; a[7]=6'd55; a[8]=6'd24; a[9]=6'd27; a[10]=6'd16; a[11]=6'd18; a[12]=6'd33; a[13]=6'd28; a[14]=6'd62; a[15]=6'd41; a[16]=6'd21; a[17]=6'd15;  end
	6'd35 : begin a[0]=6'd28; a[1]=6'd31; a[2]=6'd59; a[3]=6'd26; a[4]=6'd20; a[5]=6'd58; a[6]=6'd6; a[7]=6'd11; a[8]=6'd1; a[9]=6'd28; a[10]=6'd31; a[11]=6'd59; a[12]=6'd26; a[13]=6'd20; a[14]=6'd58; a[15]=6'd6; a[16]=6'd11; a[17]=6'd1;  end
	6'd36 : begin a[0]=6'd14; a[1]=6'd23; a[2]=6'd15; a[3]=6'd25; a[4]=6'd24; a[5]=6'd22; a[6]=6'd1; a[7]=6'd14; a[8]=6'd23; a[9]=6'd15; a[10]=6'd25; a[11]=6'd24; a[12]=6'd22; a[13]=6'd1; a[14]=6'd14; a[15]=6'd23; a[16]=6'd15; a[17]=6'd25;  end
	6'd37 : begin a[0]=6'd7; a[1]=6'd21; a[2]=6'd40; a[3]=6'd29; a[4]=6'd16; a[5]=6'd51; a[6]=6'd31; a[7]=6'd30; a[8]=6'd25; a[9]=6'd12; a[10]=6'd36; a[11]=6'd57; a[12]=6'd41; a[13]=6'd26; a[14]=6'd5; a[15]=6'd27; a[16]=6'd2; a[17]=6'd14;  end
	6'd38 : begin a[0]=6'd34; a[1]=6'd52; a[2]=6'd5; a[3]=6'd44; a[4]=6'd33; a[5]=6'd17; a[6]=6'd26; a[7]=6'd35; a[8]=6'd22; a[9]=6'd49; a[10]=6'd41; a[11]=6'd13; a[12]=6'd48; a[13]=6'd11; a[14]=6'd57; a[15]=6'd53; a[16]=6'd39; a[17]=6'd24;  end
	6'd39 : begin a[0]=6'd17; a[1]=6'd13; a[2]=6'd24; a[3]=6'd18; a[4]=6'd62; a[5]=6'd15; a[6]=6'd58; a[7]=6'd8; a[8]=6'd14; a[9]=6'd43; a[10]=6'd5; a[11]=6'd22; a[12]=6'd57; a[13]=6'd59; a[14]=6'd25; a[15]=6'd3; a[16]=6'd51; a[17]=6'd23;  end
	6'd40 : begin a[0]=6'd41; a[1]=6'd50; a[2]=6'd3; a[3]=6'd56; a[4]=6'd21; a[5]=6'd5; a[6]=6'd11; a[7]=6'd63; a[8]=6'd15; a[9]=6'd29; a[10]=6'd2; a[11]=6'd17; a[12]=6'd39; a[13]=6'd6; a[14]=6'd51; a[15]=6'd42; a[16]=6'd10; a[17]=6'd22;  end
	6'd41 : begin a[0]=6'd53; a[1]=6'd45; a[2]=6'd8; a[3]=6'd34; a[4]=6'd39; a[5]=6'd3; a[6]=6'd28; a[7]=6'd52; a[8]=6'd24; a[9]=6'd37; a[10]=6'd42; a[11]=6'd5; a[12]=6'd36; a[13]=6'd31; a[14]=6'd40; a[15]=6'd44; a[16]=6'd61; a[17]=6'd15;  end
	6'd42 : begin a[0]=6'd59; a[1]=6'd58; a[2]=6'd1; a[3]=6'd59; a[4]=6'd58; a[5]=6'd1; a[6]=6'd59; a[7]=6'd58; a[8]=6'd1; a[9]=6'd59; a[10]=6'd58; a[11]=6'd1; a[12]=6'd59; a[13]=6'd58; a[14]=6'd1; a[15]=6'd59; a[16]=6'd58; a[17]=6'd1;  end
	6'd43 : begin a[0]=6'd60; a[1]=6'd47; a[2]=6'd57; a[3]=6'd38; a[4]=6'd44; a[5]=6'd62; a[6]=6'd20; a[7]=6'd36; a[8]=6'd23; a[9]=6'd35; a[10]=6'd37; a[11]=6'd43; a[12]=6'd12; a[13]=6'd28; a[14]=6'd13; a[15]=6'd32; a[16]=6'd34; a[17]=6'd25;  end
	6'd44 : begin a[0]=6'd30; a[1]=6'd27; a[2]=6'd62; a[3]=6'd10; a[4]=6'd9; a[5]=6'd43; a[6]=6'd6; a[7]=6'd7; a[8]=6'd25; a[9]=6'd2; a[10]=6'd60; a[11]=6'd54; a[12]=6'd63; a[13]=6'd20; a[14]=6'd18; a[15]=6'd21; a[16]=6'd12; a[17]=6'd14;  end
	6'd45 : begin a[0]=6'd15; a[1]=6'd22; a[2]=6'd23; a[3]=6'd24; a[4]=6'd14; a[5]=6'd25; a[6]=6'd1; a[7]=6'd15; a[8]=6'd22; a[9]=6'd23; a[10]=6'd24; a[11]=6'd14; a[12]=6'd25; a[13]=6'd1; a[14]=6'd15; a[15]=6'd22; a[16]=6'd23; a[17]=6'd24;  end
	6'd46 : begin a[0]=6'd38; a[1]=6'd36; a[2]=6'd43; a[3]=6'd32; a[4]=6'd53; a[5]=6'd54; a[6]=6'd31; a[7]=6'd48; a[8]=6'd14; a[9]=6'd45; a[10]=6'd49; a[11]=6'd40; a[12]=6'd9; a[13]=6'd26; a[14]=6'd8; a[15]=6'd60; a[16]=6'd44; a[17]=6'd23;  end
	6'd47 : begin a[0]=6'd19; a[1]=6'd9; a[2]=6'd13; a[3]=6'd2; a[4]=6'd38; a[5]=6'd18; a[6]=6'd26; a[7]=6'd4; a[8]=6'd15; a[9]=6'd36; a[10]=6'd52; a[11]=6'd8; a[12]=6'd30; a[13]=6'd11; a[14]=6'd43; a[15]=6'd16; a[16]=6'd60; a[17]=6'd22;  end
	6'd48 : begin a[0]=6'd40; a[1]=6'd51; a[2]=6'd25; a[3]=6'd57; a[4]=6'd5; a[5]=6'd14; a[6]=6'd58; a[7]=6'd62; a[8]=6'd24; a[9]=6'd17; a[10]=6'd54; a[11]=6'd23; a[12]=6'd3; a[13]=6'd59; a[14]=6'd22; a[15]=6'd43; a[16]=6'd8; a[17]=6'd15;  end
	6'd49 : begin a[0]=6'd20; a[1]=6'd28; a[2]=6'd58; a[3]=6'd31; a[4]=6'd6; a[5]=6'd59; a[6]=6'd11; a[7]=6'd26; a[8]=6'd1; a[9]=6'd20; a[10]=6'd28; a[11]=6'd58; a[12]=6'd31; a[13]=6'd6; a[14]=6'd59; a[15]=6'd11; a[16]=6'd26; a[17]=6'd1;  end
	6'd50 : begin a[0]=6'd10; a[1]=6'd7; a[2]=6'd54; a[3]=6'd21; a[4]=6'd4; a[5]=6'd40; a[6]=6'd28; a[7]=6'd29; a[8]=6'd23; a[9]=6'd16; a[10]=6'd38; a[11]=6'd51; a[12]=6'd55; a[13]=6'd31; a[14]=6'd3; a[15]=6'd30; a[16]=6'd9; a[17]=6'd25;  end
	6'd51 : begin a[0]=6'd5; a[1]=6'd17; a[2]=6'd22; a[3]=6'd13; a[4]=6'd57; a[5]=6'd24; a[6]=6'd59; a[7]=6'd18; a[8]=6'd25; a[9]=6'd62; a[10]=6'd3; a[11]=6'd15; a[12]=6'd51; a[13]=6'd58; a[14]=6'd23; a[15]=6'd8; a[16]=6'd40; a[17]=6'd14;  end
	6'd52 : begin a[0]=6'd35; a[1]=6'd53; a[2]=6'd18; a[3]=6'd45; a[4]=6'd46; a[5]=6'd8; a[6]=6'd20; a[7]=6'd34; a[8]=6'd22; a[9]=6'd39; a[10]=6'd63; a[11]=6'd3; a[12]=6'd38; a[13]=6'd28; a[14]=6'd54; a[15]=6'd52; a[16]=6'd49; a[17]=6'd24;  end
	6'd53 : begin a[0]=6'd48; a[1]=6'd60; a[2]=6'd51; a[3]=6'd47; a[4]=6'd52; a[5]=6'd57; a[6]=6'd6; a[7]=6'd38; a[8]=6'd14; a[9]=6'd44; a[10]=6'd39; a[11]=6'd62; a[12]=6'd16; a[13]=6'd20; a[14]=6'd17; a[15]=6'd36; a[16]=6'd45; a[17]=6'd23;  end
	6'd54 : begin a[0]=6'd24; a[1]=6'd15; a[2]=6'd14; a[3]=6'd22; a[4]=6'd25; a[5]=6'd23; a[6]=6'd1; a[7]=6'd24; a[8]=6'd15; a[9]=6'd14; a[10]=6'd22; a[11]=6'd25; a[12]=6'd23; a[13]=6'd1; a[14]=6'd24; a[15]=6'd15; a[16]=6'd14; a[17]=6'd22;  end
	6'd55 : begin a[0]=6'd12; a[1]=6'd19; a[2]=6'd17; a[3]=6'd9; a[4]=6'd47; a[5]=6'd13; a[6]=6'd31; a[7]=6'd2; a[8]=6'd24; a[9]=6'd38; a[10]=6'd34; a[11]=6'd18; a[12]=6'd29; a[13]=6'd26; a[14]=6'd62; a[15]=6'd4; a[16]=6'd48; a[17]=6'd15;  end
	6'd56 : begin a[0]=6'd6; a[1]=6'd20; a[2]=6'd59; a[3]=6'd28; a[4]=6'd11; a[5]=6'd58; a[6]=6'd26; a[7]=6'd31; a[8]=6'd1; a[9]=6'd6; a[10]=6'd20; a[11]=6'd59; a[12]=6'd28; a[13]=6'd11; a[14]=6'd58; a[15]=6'd26; a[16]=6'd31; a[17]=6'd1;  end
	6'd57 : begin a[0]=6'd3; a[1]=6'd5; a[2]=6'd15; a[3]=6'd17; a[4]=6'd51; a[5]=6'd22; a[6]=6'd58; a[7]=6'd13; a[8]=6'd23; a[9]=6'd57; a[10]=6'd8; a[11]=6'd24; a[12]=6'd40; a[13]=6'd59; a[14]=6'd14; a[15]=6'd18; a[16]=6'd54; a[17]=6'd25;  end
	6'd58 : begin a[0]=6'd32; a[1]=6'd48; a[2]=6'd40; a[3]=6'd60; a[4]=6'd34; a[5]=6'd51; a[6]=6'd11; a[7]=6'd47; a[8]=6'd25; a[9]=6'd52; a[10]=6'd46; a[11]=6'd57; a[12]=6'd4; a[13]=6'd6; a[14]=6'd5; a[15]=6'd38; a[16]=6'd53; a[17]=6'd14;  end
	6'd59 : begin a[0]=6'd16; a[1]=6'd12; a[2]=6'd5; a[3]=6'd19; a[4]=6'd60; a[5]=6'd17; a[6]=6'd28; a[7]=6'd9; a[8]=6'd22; a[9]=6'd47; a[10]=6'd45; a[11]=6'd13; a[12]=6'd21; a[13]=6'd31; a[14]=6'd57; a[15]=6'd2; a[16]=6'd32; a[17]=6'd24;  end
	6'd60 : begin a[0]=6'd8; a[1]=6'd3; a[2]=6'd24; a[3]=6'd5; a[4]=6'd40; a[5]=6'd15; a[6]=6'd59; a[7]=6'd17; a[8]=6'd14; a[9]=6'd51; a[10]=6'd18; a[11]=6'd22; a[12]=6'd54; a[13]=6'd58; a[14]=6'd25; a[15]=6'd13; a[16]=6'd43; a[17]=6'd23;  end
	6'd61 : begin a[0]=6'd4; a[1]=6'd16; a[2]=6'd3; a[3]=6'd12; a[4]=6'd48; a[5]=6'd5; a[6]=6'd20; a[7]=6'd19; a[8]=6'd15; a[9]=6'd60; a[10]=6'd53; a[11]=6'd17; a[12]=6'd7; a[13]=6'd28; a[14]=6'd51; a[15]=6'd9; a[16]=6'd36; a[17]=6'd22;  end
	6'd62 : begin a[0]=6'd2; a[1]=6'd4; a[2]=6'd8; a[3]=6'd16; a[4]=6'd32; a[5]=6'd3; a[6]=6'd6; a[7]=6'd12; a[8]=6'd24; a[9]=6'd48; a[10]=6'd35; a[11]=6'd5; a[12]=6'd10; a[13]=6'd20; a[14]=6'd40; a[15]=6'd19; a[16]=6'd38; a[17]=6'd15;  end
	6'd63 : begin a[0]=6'd1; a[1]=6'd1; a[2]=6'd1; a[3]=6'd1; a[4]=6'd1; a[5]=6'd1; a[6]=6'd1; a[7]=6'd1; a[8]=6'd1; a[9]=6'd1; a[10]=6'd1; a[11]=6'd1; a[12]=6'd1; a[13]=6'd1; a[14]=6'd1; a[15]=6'd1; a[16]=6'd1; a[17]=6'd1;  end
	endcase
	return a;
endfunction



function Bit#(6) gf_inv(Bit#(6) a);
        Bit#(6) c = case(a) matches
                        6'd00 : 2;
                        6'd01 : 1;
                        6'd02 : 33;
                        6'd03 : 62;
                        6'd04 : 49;
                        6'd05 : 43;
                        6'd06 : 31;
                        6'd07 : 44;
                        6'd08 : 57;
                        6'd09 : 37;
                        6'd10 : 52;
                        6'd11 : 28;
                        6'd12 : 46;
                        6'd13 : 40;
                        6'd14 : 22;
                        6'd15 : 25;
                        6'd16 : 61;
                        6'd17 : 54;
                        6'd18 : 51;
                        6'd19 : 39;
                        6'd20 : 26;
                        6'd21 : 35;
                        6'd22 : 14;
                        6'd23 : 24;
                        6'd24 : 23;
                        6'd25 : 15;
                        6'd26 : 20;
                        6'd27 : 34;
                        6'd28 : 11;
                        6'd29 : 53;
                        6'd30 : 45;
                        6'd31 : 6;
                        6'd32 : 63;
                        6'd33 : 2;
                        6'd34 : 27;
                        6'd35 : 21;
                        6'd36 : 56;
                        6'd37 : 9;
                        6'd38 : 50;
                        6'd39 : 19;
                        6'd40 : 13;
                        6'd41 : 47;
                        6'd42 : 48;
                        6'd43 : 5;
                        6'd44 : 7;
                        6'd45 : 30;
                        6'd46 : 12;
                        6'd47 : 41;
                        6'd48 : 42;
                        6'd49 : 4;
                        6'd50 : 38;
                        6'd51 : 18;
                        6'd52 : 10;
                        6'd53 : 29;
                        6'd54 : 17;
                        6'd55 : 60;
                        6'd56 : 36;
                        6'd57 : 8;
                        6'd58 : 59;
                        6'd59 : 58;
                        6'd60 : 55;
                        6'd61 : 16;
                        6'd62 : 3;
                        6'd63 : 32;
                endcase;
        return c;
endfunction



endpackage: RS_common

