import Vector::*;

(* noinline *)
function Bit#(300) update_g(Bit#(300) g, Bit#(64) r);
	Bit#(300) g_next;
	g_next[0] = r[63]^r[48]^r[34]^r[33]^r[20]^r[18]^r[6]^r[5]^r[4]^r[3]^g[7]^g[11];
	g_next[1] = r[62]^r[48]^r[47]^r[34]^r[32]^r[20]^r[19]^r[18]^r[17]^r[6]^r[2]^g[7]^g[8]^g[11]^g[12];
	g_next[2] = r[61]^r[47]^r[46]^r[33]^r[31]^r[19]^r[18]^r[17]^r[16]^r[5]^r[1]^g[8]^g[9]^g[12]^g[13];
	g_next[3] = r[60]^r[46]^r[45]^r[32]^r[30]^r[18]^r[17]^r[16]^r[15]^r[4]^r[0]^g[9]^g[10]^g[13]^g[14];
	g_next[4] = r[59]^r[45]^r[44]^r[31]^r[29]^r[17]^r[16]^r[15]^r[14]^r[3]^g[0]^g[10]^g[11]^g[14];
	g_next[5] = r[58]^r[44]^r[43]^r[30]^r[28]^r[16]^r[15]^r[14]^r[13]^r[2]^g[1]^g[11]^g[12];
	g_next[6] = r[57]^r[43]^r[42]^r[29]^r[27]^r[15]^r[14]^r[13]^r[12]^r[1]^g[2]^g[12]^g[13];
	g_next[7] = r[56]^r[42]^r[41]^r[28]^r[26]^r[14]^r[13]^r[12]^r[11]^r[0]^g[3]^g[13]^g[14];
	g_next[8] = r[55]^r[41]^r[40]^r[27]^r[25]^r[13]^r[12]^r[11]^r[10]^g[0]^g[4]^g[14];
	g_next[9] = r[54]^r[40]^r[39]^r[26]^r[24]^r[12]^r[11]^r[10]^r[9]^g[1]^g[5];
	g_next[10] = r[53]^r[39]^r[38]^r[25]^r[23]^r[11]^r[10]^r[9]^r[8]^g[2]^g[6];
	g_next[11] = r[52]^r[38]^r[37]^r[24]^r[22]^r[10]^r[9]^r[8]^r[7]^g[3]^g[7];
	g_next[12] = r[51]^r[37]^r[36]^r[23]^r[21]^r[9]^r[8]^r[7]^r[6]^g[4]^g[8];
	g_next[13] = r[50]^r[36]^r[35]^r[22]^r[20]^r[8]^r[7]^r[6]^r[5]^g[5]^g[9];
	g_next[14] = r[49]^r[35]^r[34]^r[21]^r[19]^r[7]^r[6]^r[5]^r[4]^g[6]^g[10];
	g_next[15] = r[63]^r[58]^r[53]^r[48]^r[44]^r[43]^r[38]^r[33]^r[30]^r[28]^r[25]^r[24]^r[23]^r[18]^r[16]^r[13]^r[8]^r[6]^r[4]^r[3]^r[2]^g[18]^g[20]^g[21]^g[24]^g[25]^g[28]^g[29];
	g_next[16] = r[58]^r[48]^r[44]^r[39]^r[38]^r[34]^r[30]^r[29]^r[28]^r[18]^r[16]^r[11]^r[8]^r[4]^r[2]^g[15]^g[18]^g[19]^g[20]^g[22]^g[24]^g[26]^g[28];
	g_next[17] = r[53]^r[48]^r[39]^r[33]^r[29]^r[28]^r[25]^r[20]^r[15]^r[13]^r[11]^r[10]^r[8]^r[5]^r[0]^g[15]^g[16]^g[19]^g[20]^g[21]^g[23]^g[25]^g[27]^g[29];
	g_next[18] = r[62]^r[57]^r[52]^r[48]^r[47]^r[42]^r[37]^r[34]^r[32]^r[29]^r[28]^r[27]^r[22]^r[20]^r[17]^r[12]^r[10]^r[8]^r[7]^r[6]^r[2]^r[1]^r[0]^g[16]^g[17]^g[20]^g[21]^g[22]^g[24]^g[26]^g[28];
	g_next[19] = r[57]^r[47]^r[43]^r[38]^r[37]^r[33]^r[29]^r[28]^r[27]^r[17]^r[15]^r[10]^r[7]^r[3]^r[1]^g[17]^g[18]^g[21]^g[22]^g[23]^g[25]^g[27]^g[29];
	g_next[20] = r[52]^r[47]^r[38]^r[32]^r[28]^r[27]^r[24]^r[19]^r[14]^r[12]^r[10]^r[9]^r[7]^r[4]^g[15]^g[18]^g[19]^g[22]^g[23]^g[24]^g[26]^g[28];
	g_next[21] = r[61]^r[56]^r[51]^r[47]^r[46]^r[41]^r[36]^r[33]^r[31]^r[28]^r[27]^r[26]^r[21]^r[19]^r[16]^r[11]^r[9]^r[7]^r[6]^r[5]^r[1]^r[0]^g[15]^g[16]^g[19]^g[20]^g[23]^g[24]^g[25]^g[27]^g[29];
	g_next[22] = r[56]^r[46]^r[42]^r[37]^r[36]^r[32]^r[28]^r[27]^r[26]^r[16]^r[14]^r[9]^r[6]^r[2]^r[0]^g[16]^g[17]^g[20]^g[21]^g[24]^g[25]^g[26]^g[28];
	g_next[23] = r[51]^r[46]^r[37]^r[31]^r[27]^r[26]^r[23]^r[18]^r[13]^r[11]^r[9]^r[8]^r[6]^r[3]^g[17]^g[18]^g[21]^g[22]^g[25]^g[26]^g[27]^g[29];
	g_next[24] = r[60]^r[55]^r[50]^r[46]^r[45]^r[40]^r[35]^r[32]^r[30]^r[27]^r[26]^r[25]^r[20]^r[18]^r[15]^r[10]^r[8]^r[6]^r[5]^r[4]^r[0]^g[15]^g[18]^g[19]^g[22]^g[23]^g[26]^g[27]^g[28];
	g_next[25] = r[55]^r[45]^r[41]^r[36]^r[35]^r[31]^r[27]^r[26]^r[25]^r[15]^r[13]^r[8]^r[5]^r[1]^g[15]^g[16]^g[19]^g[20]^g[23]^g[24]^g[27]^g[28]^g[29];
	g_next[26] = r[50]^r[45]^r[36]^r[30]^r[26]^r[25]^r[22]^r[17]^r[12]^r[10]^r[8]^r[7]^r[5]^r[2]^g[16]^g[17]^g[20]^g[21]^g[24]^g[25]^g[28]^g[29];
	g_next[27] = r[59]^r[54]^r[49]^r[45]^r[44]^r[39]^r[34]^r[31]^r[29]^r[26]^r[25]^r[24]^r[19]^r[17]^r[14]^r[9]^r[7]^r[5]^r[4]^r[3]^g[15]^g[17]^g[18]^g[21]^g[22]^g[25]^g[26]^g[29];
	g_next[28] = r[54]^r[44]^r[40]^r[35]^r[34]^r[30]^r[26]^r[25]^r[24]^r[14]^r[12]^r[7]^r[4]^r[0]^g[16]^g[18]^g[19]^g[22]^g[23]^g[26]^g[27];
	g_next[29] = r[49]^r[44]^r[35]^r[29]^r[25]^r[24]^r[21]^r[16]^r[11]^r[9]^r[7]^r[6]^r[4]^r[1]^g[17]^g[19]^g[20]^g[23]^g[24]^g[27]^g[28];
	g_next[30] = r[63]^r[60]^r[57]^r[54]^r[51]^r[48]^r[46]^r[45]^r[42]^r[40]^r[39]^r[36]^r[33]^r[32]^r[30]^r[29]^r[27]^r[24]^r[22]^r[21]^r[20]^r[17]^r[16]^r[15]^r[12]^r[9]^r[6]^r[4]^r[3]^r[1]^r[0]^g[33]^g[36]^g[37]^g[40];
	g_next[31] = r[60]^r[54]^r[48]^r[46]^r[43]^r[42]^r[36]^r[32]^r[30]^r[24]^r[22]^r[20]^r[19]^r[15]^r[9]^r[4]^r[3]^g[33]^g[34]^g[36]^g[38]^g[40]^g[41];
	g_next[32] = r[57]^r[54]^r[45]^r[43]^r[42]^r[33]^r[30]^r[29]^r[26]^r[23]^r[21]^r[20]^r[19]^r[18]^r[15]^r[6]^r[3]^r[1]^g[34]^g[35]^g[37]^g[39]^g[41]^g[42];
	g_next[33] = r[54]^r[42]^r[40]^r[37]^r[34]^r[31]^r[30]^r[28]^r[26]^r[25]^r[22]^r[20]^r[19]^r[18]^r[12]^r[9]^r[6]^r[0]^g[35]^g[36]^g[38]^g[40]^g[42]^g[43];
	g_next[34] = r[51]^r[48]^r[45]^r[42]^r[37]^r[31]^r[27]^r[25]^r[24]^r[23]^r[21]^r[20]^r[19]^r[18]^r[9]^r[3]^r[0]^g[36]^g[37]^g[39]^g[41]^g[43]^g[44];
	g_next[35] = r[62]^r[59]^r[56]^r[53]^r[50]^r[48]^r[47]^r[44]^r[42]^r[41]^r[38]^r[35]^r[34]^r[32]^r[31]^r[29]^r[26]^r[24]^r[23]^r[22]^r[19]^r[18]^r[17]^r[14]^r[11]^r[8]^r[6]^r[5]^r[3]^r[2]^g[30]^g[37]^g[38]^g[40]^g[42]^g[44];
	g_next[36] = r[59]^r[53]^r[47]^r[45]^r[42]^r[41]^r[35]^r[31]^r[29]^r[23]^r[21]^r[19]^r[18]^r[14]^r[8]^r[3]^r[2]^g[31]^g[38]^g[39]^g[41]^g[43];
	g_next[37] = r[56]^r[53]^r[44]^r[42]^r[41]^r[32]^r[29]^r[28]^r[25]^r[22]^r[20]^r[19]^r[18]^r[17]^r[14]^r[5]^r[2]^r[0]^g[32]^g[39]^g[40]^g[42]^g[44];
	g_next[38] = r[53]^r[41]^r[39]^r[36]^r[33]^r[30]^r[29]^r[27]^r[25]^r[24]^r[21]^r[19]^r[18]^r[17]^r[11]^r[8]^r[5]^g[30]^g[33]^g[40]^g[41]^g[43];
	g_next[39] = r[50]^r[47]^r[44]^r[41]^r[36]^r[30]^r[26]^r[24]^r[23]^r[22]^r[20]^r[19]^r[18]^r[17]^r[8]^r[2]^g[30]^g[31]^g[34]^g[41]^g[42]^g[44];
	g_next[40] = r[61]^r[58]^r[55]^r[52]^r[49]^r[47]^r[46]^r[43]^r[41]^r[40]^r[37]^r[34]^r[33]^r[31]^r[30]^r[28]^r[25]^r[23]^r[22]^r[21]^r[18]^r[17]^r[16]^r[13]^r[10]^r[7]^r[5]^r[4]^r[2]^r[1]^g[31]^g[32]^g[35]^g[42]^g[43];
	g_next[41] = r[58]^r[52]^r[46]^r[44]^r[41]^r[40]^r[34]^r[30]^r[28]^r[22]^r[20]^r[18]^r[17]^r[13]^r[7]^r[2]^r[1]^g[32]^g[33]^g[36]^g[43]^g[44];
	g_next[42] = r[55]^r[52]^r[43]^r[41]^r[40]^r[31]^r[28]^r[27]^r[24]^r[21]^r[19]^r[18]^r[17]^r[16]^r[13]^r[4]^r[1]^g[30]^g[33]^g[34]^g[37]^g[44];
	g_next[43] = r[52]^r[40]^r[38]^r[35]^r[32]^r[29]^r[28]^r[26]^r[24]^r[23]^r[20]^r[18]^r[17]^r[16]^r[10]^r[7]^r[4]^g[31]^g[34]^g[35]^g[38];
	g_next[44] = r[49]^r[46]^r[43]^r[40]^r[35]^r[29]^r[25]^r[23]^r[22]^r[21]^r[19]^r[18]^r[17]^r[16]^r[7]^r[1]^g[32]^g[35]^g[36]^g[39];
	g_next[45] = r[63]^r[48]^r[46]^r[33]^r[32]^r[30]^r[29]^r[18]^r[12]^r[3]^r[2]^r[1]^g[46]^g[49]^g[51]^g[53]^g[55]^g[57]^g[59];
	g_next[46] = r[50]^r[48]^r[35]^r[34]^r[32]^r[31]^r[20]^r[14]^r[5]^r[4]^r[3]^g[45]^g[46]^g[47]^g[49]^g[50]^g[51]^g[52]^g[53]^g[54]^g[55]^g[56]^g[57]^g[58]^g[59];
	g_next[47] = r[52]^r[48]^r[37]^r[36]^r[35]^r[33]^r[32]^r[31]^r[22]^r[20]^r[16]^r[14]^r[7]^r[6]^r[4]^r[3]^r[1]^r[0]^g[46]^g[47]^g[48]^g[50]^g[51]^g[52]^g[53]^g[54]^g[55]^g[56]^g[57]^g[58]^g[59];
	g_next[48] = r[54]^r[52]^r[50]^r[48]^r[39]^r[38]^r[36]^r[34]^r[32]^r[31]^r[24]^r[20]^r[18]^r[14]^r[9]^r[8]^r[7]^r[5]^r[4]^r[2]^r[1]^g[45]^g[47]^g[48]^g[49]^g[51]^g[52]^g[53]^g[54]^g[55]^g[56]^g[57]^g[58]^g[59];
	g_next[49] = r[56]^r[48]^r[41]^r[40]^r[39]^r[33]^r[32]^r[31]^r[26]^r[24]^r[22]^r[18]^r[16]^r[14]^r[11]^r[10]^r[8]^r[6]^r[5]^r[3]^r[2]^r[0]^g[46]^g[48]^g[49]^g[50]^g[52]^g[53]^g[54]^g[55]^g[56]^g[57]^g[58]^g[59];
	g_next[50] = r[58]^r[56]^r[50]^r[48]^r[43]^r[42]^r[40]^r[39]^r[35]^r[34]^r[32]^r[31]^r[28]^r[22]^r[20]^r[14]^r[13]^r[12]^r[11]^r[7]^r[6]^r[4]^r[3]^g[45]^g[47]^g[49]^g[50]^g[51]^g[53]^g[54]^g[55]^g[56]^g[57]^g[58]^g[59];
	g_next[51] = r[60]^r[56]^r[52]^r[48]^r[45]^r[44]^r[43]^r[41]^r[40]^r[39]^r[37]^r[36]^r[35]^r[33]^r[32]^r[31]^r[30]^r[28]^r[24]^r[20]^r[16]^r[15]^r[12]^r[11]^r[9]^r[8]^r[7]^r[5]^r[4]^r[3]^r[1]^g[46]^g[48]^g[50]^g[51]^g[52]^g[54]^g[55]^g[56]^g[57]^g[58]^g[59];
	g_next[52] = r[62]^r[60]^r[58]^r[56]^r[54]^r[52]^r[50]^r[48]^r[47]^r[46]^r[44]^r[42]^r[40]^r[38]^r[36]^r[34]^r[31]^r[28]^r[26]^r[24]^r[22]^r[20]^r[18]^r[17]^r[16]^r[15]^r[14]^r[13]^r[12]^r[10]^r[8]^r[6]^r[4]^r[1]^r[0]^g[45]^g[47]^g[49]^g[51]^g[52]^g[53]^g[55]^g[56]^g[57]^g[58]^g[59];
	g_next[53] = r[49]^r[47]^r[34]^r[33]^r[31]^r[30]^r[19]^r[13]^r[4]^r[3]^r[2]^g[46]^g[48]^g[50]^g[52]^g[53]^g[54]^g[56]^g[57]^g[58]^g[59];
	g_next[54] = r[51]^r[47]^r[36]^r[35]^r[34]^r[32]^r[31]^r[30]^r[21]^r[19]^r[15]^r[13]^r[6]^r[5]^r[3]^r[2]^r[0]^g[45]^g[47]^g[49]^g[51]^g[53]^g[54]^g[55]^g[57]^g[58]^g[59];
	g_next[55] = r[53]^r[51]^r[49]^r[47]^r[38]^r[37]^r[35]^r[33]^r[31]^r[30]^r[23]^r[19]^r[17]^r[13]^r[8]^r[7]^r[6]^r[4]^r[3]^r[1]^r[0]^g[46]^g[48]^g[50]^g[52]^g[54]^g[55]^g[56]^g[58]^g[59];
	g_next[56] = r[55]^r[47]^r[40]^r[39]^r[38]^r[32]^r[31]^r[30]^r[25]^r[23]^r[21]^r[17]^r[15]^r[13]^r[10]^r[9]^r[7]^r[5]^r[4]^r[2]^r[1]^g[45]^g[47]^g[49]^g[51]^g[53]^g[55]^g[56]^g[57]^g[59];
	g_next[57] = r[57]^r[55]^r[49]^r[47]^r[42]^r[41]^r[39]^r[38]^r[34]^r[33]^r[31]^r[30]^r[27]^r[21]^r[19]^r[13]^r[12]^r[11]^r[10]^r[6]^r[5]^r[3]^r[2]^g[46]^g[48]^g[50]^g[52]^g[54]^g[56]^g[57]^g[58];
	g_next[58] = r[59]^r[55]^r[51]^r[47]^r[44]^r[43]^r[42]^r[40]^r[39]^r[38]^r[36]^r[35]^r[34]^r[32]^r[31]^r[30]^r[29]^r[27]^r[23]^r[19]^r[15]^r[14]^r[11]^r[10]^r[8]^r[7]^r[6]^r[4]^r[3]^r[2]^r[0]^g[47]^g[49]^g[51]^g[53]^g[55]^g[57]^g[58]^g[59];
	g_next[59] = r[61]^r[59]^r[57]^r[55]^r[53]^r[51]^r[49]^r[47]^r[46]^r[45]^r[43]^r[41]^r[39]^r[37]^r[35]^r[33]^r[30]^r[27]^r[25]^r[23]^r[21]^r[19]^r[17]^r[16]^r[15]^r[14]^r[13]^r[12]^r[11]^r[9]^r[7]^r[5]^r[3]^r[0]^g[45]^g[48]^g[50]^g[52]^g[54]^g[56]^g[58]^g[59];
	g_next[60] = r[63]^r[58]^r[53]^r[52]^r[50]^r[48]^r[44]^r[43]^r[41]^r[37]^r[33]^r[30]^r[28]^r[25]^r[24]^r[23]^r[20]^r[19]^r[18]^r[16]^r[11]^r[8]^r[3]^r[2]^r[0]^g[63]^g[65]^g[69]^g[73]^g[74];
	g_next[61] = r[58]^r[55]^r[52]^r[48]^r[40]^r[39]^r[33]^r[30]^r[27]^r[25]^r[24]^r[23]^r[20]^r[19]^r[15]^r[13]^r[12]^r[10]^r[8]^r[2]^r[0]^g[60]^g[63]^g[64]^g[65]^g[66]^g[69]^g[70]^g[73];
	g_next[62] = r[58]^r[55]^r[53]^r[47]^r[42]^r[41]^r[39]^r[38]^r[30]^r[27]^r[25]^r[23]^r[22]^r[19]^r[18]^r[17]^r[14]^r[13]^r[12]^r[8]^r[3]^r[2]^g[60]^g[61]^g[64]^g[65]^g[66]^g[67]^g[70]^g[71]^g[74];
	g_next[63] = r[61]^r[58]^r[56]^r[51]^r[46]^r[44]^r[42]^r[41]^r[40]^r[39]^r[38]^r[36]^r[33]^r[31]^r[30]^r[28]^r[26]^r[25]^r[21]^r[18]^r[17]^r[13]^r[12]^r[11]^r[8]^r[6]^r[5]^r[2]^r[1]^r[0]^g[61]^g[62]^g[65]^g[66]^g[67]^g[68]^g[71]^g[72];
	g_next[64] = r[61]^r[53]^r[51]^r[47]^r[43]^r[41]^r[39]^r[38]^r[36]^r[33]^r[28]^r[26]^r[25]^r[19]^r[17]^r[16]^r[15]^r[14]^r[12]^r[11]^r[8]^r[5]^r[1]^g[62]^g[63]^g[66]^g[67]^g[68]^g[69]^g[72]^g[73];
	g_next[65] = r[51]^r[50]^r[46]^r[45]^r[40]^r[39]^r[38]^r[36]^r[31]^r[22]^r[20]^r[18]^r[16]^r[15]^r[13]^r[12]^r[8]^r[1]^g[63]^g[64]^g[67]^g[68]^g[69]^g[70]^g[73]^g[74];
	g_next[66] = r[59]^r[54]^r[53]^r[51]^r[49]^r[45]^r[44]^r[42]^r[38]^r[34]^r[31]^r[29]^r[26]^r[25]^r[24]^r[21]^r[20]^r[19]^r[17]^r[12]^r[9]^r[4]^r[3]^r[1]^g[60]^g[64]^g[65]^g[68]^g[69]^g[70]^g[71]^g[74];
	g_next[67] = r[56]^r[54]^r[51]^r[45]^r[44]^r[42]^r[41]^r[40]^r[38]^r[29]^r[28]^r[19]^r[17]^r[16]^r[14]^r[13]^r[12]^r[11]^r[4]^r[0]^g[61]^g[65]^g[66]^g[69]^g[70]^g[71]^g[72];
	g_next[68] = r[59]^r[51]^r[48]^r[45]^r[44]^r[43]^r[41]^r[39]^r[38]^r[31]^r[29]^r[26]^r[24]^r[23]^r[20]^r[18]^r[17]^r[16]^r[15]^r[12]^r[11]^r[9]^r[3]^g[62]^g[66]^g[67]^g[70]^g[71]^g[72]^g[73];
	g_next[69] = r[62]^r[57]^r[52]^r[51]^r[48]^r[47]^r[44]^r[42]^r[40]^r[38]^r[37]^r[34]^r[32]^r[27]^r[24]^r[23]^r[22]^r[20]^r[19]^r[17]^r[16]^r[15]^r[14]^r[13]^r[11]^r[7]^r[6]^r[2]^r[1]^g[63]^g[67]^g[68]^g[71]^g[72]^g[73]^g[74];
	g_next[70] = r[57]^r[54]^r[51]^r[47]^r[39]^r[38]^r[32]^r[29]^r[26]^r[24]^r[23]^r[22]^r[19]^r[18]^r[14]^r[12]^r[11]^r[9]^r[7]^r[1]^g[60]^g[64]^g[68]^g[69]^g[72]^g[73]^g[74];
	g_next[71] = r[57]^r[54]^r[52]^r[46]^r[41]^r[40]^r[38]^r[37]^r[29]^r[26]^r[24]^r[22]^r[21]^r[18]^r[17]^r[16]^r[13]^r[12]^r[11]^r[7]^r[2]^r[1]^g[61]^g[65]^g[69]^g[70]^g[73]^g[74];
	g_next[72] = r[60]^r[57]^r[55]^r[50]^r[45]^r[43]^r[41]^r[40]^r[39]^r[38]^r[37]^r[35]^r[32]^r[30]^r[29]^r[27]^r[25]^r[24]^r[20]^r[17]^r[16]^r[12]^r[11]^r[10]^r[7]^r[5]^r[4]^r[1]^r[0]^g[60]^g[62]^g[66]^g[70]^g[71]^g[74];
	g_next[73] = r[60]^r[52]^r[50]^r[46]^r[42]^r[40]^r[38]^r[37]^r[35]^r[32]^r[27]^r[25]^r[24]^r[18]^r[16]^r[15]^r[14]^r[13]^r[11]^r[10]^r[7]^r[4]^r[0]^g[61]^g[63]^g[67]^g[71]^g[72];
	g_next[74] = r[50]^r[49]^r[45]^r[44]^r[39]^r[38]^r[37]^r[35]^r[30]^r[21]^r[19]^r[17]^r[15]^r[14]^r[12]^r[11]^r[7]^r[0]^g[62]^g[64]^g[68]^g[72]^g[73];
	g_next[75] = r[63]^r[54]^r[48]^r[46]^r[45]^r[44]^r[42]^r[40]^r[36]^r[33]^r[29]^r[27]^r[26]^r[25]^r[24]^r[21]^r[20]^r[18]^r[17]^r[14]^r[12]^r[9]^r[8]^r[6]^r[3]^r[0]^g[77]^g[78]^g[79]^g[80]^g[81]^g[82]^g[83]^g[84]^g[85]^g[87]^g[88];
	g_next[76] = r[59]^r[54]^r[52]^r[50]^r[48]^r[46]^r[44]^r[43]^r[40]^r[37]^r[36]^r[33]^r[32]^r[31]^r[27]^r[26]^r[24]^r[23]^r[21]^r[18]^r[14]^r[13]^r[12]^r[8]^r[7]^r[5]^r[3]^r[0]^g[77]^g[86]^g[87]^g[89];
	g_next[77] = r[59]^r[56]^r[55]^r[48]^r[45]^r[43]^r[41]^r[36]^r[32]^r[31]^r[29]^r[27]^r[26]^r[25]^r[24]^r[22]^r[21]^r[18]^r[17]^r[13]^r[11]^r[10]^r[9]^r[8]^r[7]^r[5]^r[2]^r[1]^r[0]^g[75]^g[78]^g[87]^g[88];
	g_next[78] = r[60]^r[56]^r[50]^r[48]^r[45]^r[44]^r[43]^r[41]^r[37]^r[36]^r[33]^r[32]^r[30]^r[28]^r[25]^r[23]^r[22]^r[21]^r[18]^r[15]^r[13]^r[10]^r[8]^r[7]^r[6]^r[4]^r[2]^g[75]^g[76]^g[79]^g[88]^g[89];
	g_next[79] = r[55]^r[49]^r[47]^r[46]^r[45]^r[43]^r[41]^r[37]^r[34]^r[30]^r[28]^r[27]^r[26]^r[25]^r[22]^r[21]^r[19]^r[18]^r[15]^r[13]^r[10]^r[9]^r[7]^r[4]^r[1]^g[76]^g[77]^g[80]^g[89];
	g_next[80] = r[60]^r[53]^r[51]^r[46]^r[44]^r[43]^r[38]^r[33]^r[32]^r[30]^r[26]^r[24]^r[21]^r[18]^r[14]^r[10]^r[8]^r[7]^r[6]^g[75]^g[77]^g[78]^g[81];
	g_next[81] = r[57]^r[56]^r[53]^r[51]^r[49]^r[43]^r[42]^r[38]^r[37]^r[28]^r[27]^r[25]^r[24]^r[23]^r[22]^r[21]^r[19]^r[12]^r[11]^r[9]^r[7]^r[3]^r[2]^r[1]^r[0]^g[75]^g[76]^g[78]^g[79]^g[82];
	g_next[82] = r[61]^r[56]^r[53]^r[46]^r[45]^r[44]^r[43]^r[34]^r[33]^r[31]^r[29]^r[28]^r[27]^r[26]^r[25]^r[21]^r[16]^r[14]^r[12]^r[8]^r[5]^r[2]^r[1]^g[75]^g[76]^g[77]^g[79]^g[80]^g[83];
	g_next[83] = r[61]^r[53]^r[50]^r[48]^r[47]^r[45]^r[43]^r[42]^r[38]^r[35]^r[34]^r[33]^r[25]^r[23]^r[22]^r[21]^r[20]^r[19]^r[12]^r[11]^r[10]^r[1]^g[75]^g[76]^g[77]^g[78]^g[80]^g[81]^g[84];
	g_next[84] = r[54]^r[53]^r[52]^r[50]^r[48]^r[44]^r[43]^r[42]^r[39]^r[38]^r[35]^r[31]^r[27]^r[23]^r[21]^r[20]^r[15]^r[12]^r[10]^r[9]^r[8]^r[7]^r[1]^r[0]^g[75]^g[76]^g[77]^g[78]^g[79]^g[81]^g[82]^g[85];
	g_next[85] = r[58]^r[57]^r[53]^r[48]^r[42]^r[35]^r[31]^r[29]^r[28]^r[27]^r[26]^r[25]^r[24]^r[22]^r[21]^r[15]^r[13]^r[9]^r[7]^r[4]^r[3]^r[2]^g[75]^g[76]^g[77]^g[78]^g[79]^g[80]^g[82]^g[83]^g[86];
	g_next[86] = r[62]^r[58]^r[54]^r[53]^r[48]^r[47]^r[46]^r[45]^r[44]^r[42]^r[34]^r[32]^r[31]^r[30]^r[25]^r[24]^r[21]^r[17]^r[7]^r[6]^r[4]^r[0]^g[75]^g[76]^g[77]^g[78]^g[79]^g[80]^g[81]^g[83]^g[84]^g[87];
	g_next[87] = r[58]^r[53]^r[51]^r[49]^r[47]^r[45]^r[43]^r[42]^r[39]^r[36]^r[35]^r[32]^r[31]^r[30]^r[26]^r[25]^r[23]^r[22]^r[20]^r[17]^r[13]^r[12]^r[11]^r[7]^r[6]^r[4]^r[2]^g[75]^g[76]^g[77]^g[78]^g[79]^g[80]^g[81]^g[82]^g[84]^g[85]^g[88];
	g_next[88] = r[58]^r[55]^r[54]^r[47]^r[44]^r[42]^r[40]^r[35]^r[31]^r[30]^r[28]^r[26]^r[25]^r[24]^r[23]^r[21]^r[20]^r[17]^r[16]^r[12]^r[10]^r[9]^r[8]^r[7]^r[6]^r[4]^r[1]^r[0]^g[75]^g[76]^g[77]^g[78]^g[79]^g[80]^g[81]^g[82]^g[83]^g[85]^g[86]^g[89];
	g_next[89] = r[59]^r[55]^r[49]^r[47]^r[44]^r[43]^r[42]^r[40]^r[36]^r[35]^r[32]^r[31]^r[29]^r[27]^r[24]^r[22]^r[21]^r[20]^r[17]^r[14]^r[12]^r[9]^r[7]^r[6]^r[5]^r[3]^r[1]^g[76]^g[77]^g[78]^g[79]^g[80]^g[81]^g[82]^g[83]^g[84]^g[86]^g[87];
	g_next[90] = r[63]^r[54]^r[50]^r[48]^r[46]^r[45]^r[37]^r[36]^r[33]^r[30]^r[29]^r[27]^r[24]^r[22]^r[18]^r[16]^r[14]^r[11]^r[10]^r[9]^r[3]^g[91]^g[92]^g[94]^g[95]^g[98]^g[99]^g[100]^g[102]^g[104];
	g_next[91] = r[56]^r[55]^r[52]^r[51]^r[50]^r[48]^r[46]^r[41]^r[40]^r[39]^r[36]^r[33]^r[32]^r[31]^r[30]^r[29]^r[28]^r[26]^r[25]^r[23]^r[22]^r[18]^r[16]^r[14]^r[11]^r[9]^r[8]^r[3]^r[2]^r[1]^r[0]^g[90]^g[91]^g[93]^g[94]^g[96]^g[98]^g[101]^g[102]^g[103]^g[104];
	g_next[92] = r[55]^r[51]^r[49]^r[47]^r[46]^r[38]^r[37]^r[34]^r[31]^r[30]^r[28]^r[25]^r[23]^r[19]^r[17]^r[15]^r[12]^r[11]^r[10]^r[4]^g[91]^g[92]^g[94]^g[95]^g[97]^g[99]^g[102]^g[103]^g[104];
	g_next[93] = r[57]^r[56]^r[55]^r[53]^r[52]^r[46]^r[42]^r[41]^r[40]^r[38]^r[33]^r[32]^r[29]^r[28]^r[27]^r[26]^r[25]^r[24]^r[11]^r[9]^r[3]^r[2]^r[1]^r[0]^g[90]^g[92]^g[93]^g[95]^g[96]^g[98]^g[100]^g[103]^g[104];
	g_next[94] = r[57]^r[55]^r[53]^r[50]^r[48]^r[47]^r[46]^r[42]^r[41]^r[40]^r[39]^r[35]^r[33]^r[31]^r[28]^r[27]^r[25]^r[20]^r[18]^r[16]^r[13]^r[12]^r[9]^r[5]^r[3]^r[2]^r[1]^r[0]^g[91]^g[93]^g[94]^g[96]^g[97]^g[99]^g[101]^g[104];
	g_next[95] = r[58]^r[56]^r[55]^r[54]^r[50]^r[48]^r[46]^r[43]^r[40]^r[35]^r[34]^r[31]^r[30]^r[29]^r[26]^r[20]^r[18]^r[16]^r[13]^r[10]^r[9]^r[5]^r[4]^g[90]^g[92]^g[94]^g[95]^g[97]^g[98]^g[100]^g[102];
	g_next[96] = r[55]^r[51]^r[50]^r[49]^r[47]^r[46]^r[42]^r[41]^r[36]^r[35]^r[32]^r[31]^r[30]^r[28]^r[21]^r[20]^r[19]^r[18]^r[17]^r[16]^r[14]^r[9]^r[6]^r[5]^r[3]^r[2]^r[1]^g[90]^g[91]^g[93]^g[95]^g[96]^g[98]^g[99]^g[101]^g[103];
	g_next[97] = r[59]^r[57]^r[56]^r[50]^r[46]^r[44]^r[42]^r[28]^r[27]^r[20]^r[18]^r[16]^r[11]^r[10]^r[9]^r[3]^r[2]^r[1]^r[0]^g[90]^g[91]^g[92]^g[94]^g[96]^g[97]^g[99]^g[100]^g[102]^g[104];
	g_next[98] = r[59]^r[57]^r[52]^r[51]^r[48]^r[47]^r[46]^r[44]^r[43]^r[37]^r[36]^r[33]^r[32]^r[31]^r[29]^r[28]^r[27]^r[22]^r[21]^r[19]^r[17]^r[16]^r[15]^r[11]^r[9]^r[7]^r[6]^r[4]^r[1]^g[91]^g[92]^g[93]^g[95]^g[97]^g[98]^g[100]^g[101]^g[103];
	g_next[99] = r[60]^r[59]^r[58]^r[52]^r[48]^r[46]^r[45]^r[44]^r[37]^r[36]^r[33]^r[32]^r[31]^r[27]^r[22]^r[16]^r[15]^r[12]^r[10]^r[9]^r[7]^r[6]^r[3]^r[2]^r[0]^g[92]^g[93]^g[94]^g[96]^g[98]^g[99]^g[101]^g[102]^g[104];
	g_next[100] = r[59]^r[53]^r[49]^r[47]^r[46]^r[38]^r[36]^r[34]^r[31]^r[30]^r[29]^r[28]^r[27]^r[23]^r[20]^r[18]^r[17]^r[15]^r[9]^r[8]^r[6]^r[5]^r[3]^r[0]^g[90]^g[93]^g[94]^g[95]^g[97]^g[99]^g[100]^g[102]^g[103];
	g_next[101] = r[61]^r[60]^r[45]^r[37]^r[36]^r[33]^r[32]^r[31]^r[30]^r[29]^r[27]^r[20]^r[18]^r[16]^r[15]^r[13]^r[11]^r[10]^r[9]^r[7]^r[6]^r[5]^r[4]^r[1]^r[0]^g[90]^g[91]^g[94]^g[95]^g[96]^g[98]^g[100]^g[101]^g[103]^g[104];
	g_next[102] = r[61]^r[54]^r[50]^r[48]^r[47]^r[45]^r[39]^r[36]^r[35]^r[33]^r[28]^r[27]^r[24]^r[21]^r[20]^r[19]^r[15]^r[13]^r[11]^r[5]^g[91]^g[92]^g[95]^g[96]^g[97]^g[99]^g[101]^g[102]^g[104];
	g_next[103] = r[62]^r[54]^r[50]^r[48]^r[47]^r[46]^r[45]^r[39]^r[38]^r[37]^r[36]^r[35]^r[34]^r[32]^r[31]^r[30]^r[27]^r[24]^r[20]^r[17]^r[16]^r[15]^r[14]^r[13]^r[12]^r[10]^r[8]^r[7]^r[6]^r[2]^r[1]^r[0]^g[90]^g[92]^g[93]^g[96]^g[97]^g[98]^g[100]^g[102]^g[103];
	g_next[104] = r[55]^r[54]^r[51]^r[50]^r[49]^r[47]^r[45]^r[40]^r[39]^r[38]^r[35]^r[32]^r[31]^r[30]^r[29]^r[28]^r[27]^r[25]^r[24]^r[22]^r[21]^r[17]^r[15]^r[13]^r[10]^r[8]^r[7]^r[2]^r[1]^r[0]^g[90]^g[91]^g[93]^g[94]^g[97]^g[98]^g[99]^g[101]^g[103]^g[104];
	g_next[105] = r[63]^r[62]^r[61]^r[60]^r[59]^r[58]^r[57]^r[56]^r[55]^r[54]^r[53]^r[52]^r[51]^r[50]^r[49]^r[47]^r[46]^r[45]^r[44]^r[43]^r[42]^r[41]^r[40]^r[39]^r[38]^r[37]^r[36]^r[35]^r[31]^r[30]^r[29]^r[28]^r[27]^r[26]^r[25]^r[24]^r[23]^r[22]^r[21]^r[19]^r[17]^r[15]^r[14]^r[13]^r[12]^r[11]^r[10]^r[9]^r[8]^r[7]^r[4]^r[2]^g[105]^g[112]^g[116];
	g_next[106] = r[62]^r[60]^r[58]^r[56]^r[54]^r[52]^r[50]^r[47]^r[45]^r[43]^r[41]^r[39]^r[37]^r[35]^r[34]^r[33]^r[32]^r[30]^r[28]^r[26]^r[24]^r[22]^r[19]^r[18]^r[15]^r[13]^r[11]^r[9]^r[7]^r[6]^r[5]^r[2]^r[1]^r[0]^g[106]^g[112]^g[113]^g[116]^g[117];
	g_next[107] = r[61]^r[60]^r[57]^r[56]^r[53]^r[52]^r[49]^r[48]^r[47]^r[44]^r[43]^r[40]^r[39]^r[36]^r[35]^r[33]^r[31]^r[30]^r[27]^r[26]^r[23]^r[22]^r[18]^r[14]^r[13]^r[10]^r[9]^r[6]^r[4]^r[3]^r[2]^r[0]^g[107]^g[113]^g[114]^g[117]^g[118];
	g_next[108] = r[60]^r[56]^r[52]^r[48]^r[46]^r[45]^r[44]^r[42]^r[41]^r[40]^r[38]^r[37]^r[36]^r[34]^r[33]^r[30]^r[26]^r[22]^r[17]^r[16]^r[15]^r[14]^r[12]^r[11]^r[10]^r[8]^r[7]^r[6]^r[3]^r[1]^r[0]^g[108]^g[114]^g[115]^g[118]^g[119];
	g_next[109] = r[59]^r[58]^r[57]^r[56]^r[51]^r[50]^r[49]^r[48]^r[45]^r[43]^r[42]^r[40]^r[37]^r[35]^r[34]^r[32]^r[31]^r[30]^r[25]^r[24]^r[23]^r[22]^r[16]^r[14]^r[11]^r[9]^r[8]^r[6]^r[2]^r[1]^g[105]^g[109]^g[115]^g[116]^g[119];
	g_next[110] = r[58]^r[56]^r[50]^r[48]^r[44]^r[43]^r[41]^r[40]^r[36]^r[35]^r[33]^r[32]^r[30]^r[24]^r[22]^r[15]^r[14]^r[10]^r[9]^r[7]^r[6]^r[1]^g[106]^g[110]^g[116]^g[117];
	g_next[111] = r[57]^r[56]^r[49]^r[48]^r[43]^r[40]^r[35]^r[32]^r[29]^r[28]^r[27]^r[26]^r[25]^r[24]^r[21]^r[20]^r[19]^r[18]^r[17]^r[16]^r[15]^r[13]^r[12]^r[11]^r[10]^r[8]^r[7]^r[5]^r[4]^r[3]^r[2]^r[1]^g[107]^g[111]^g[117]^g[118];
	g_next[112] = r[56]^r[48]^r[42]^r[41]^r[40]^r[34]^r[33]^r[32]^r[28]^r[26]^r[24]^r[20]^r[18]^r[16]^r[14]^r[13]^r[11]^r[9]^r[8]^r[6]^r[5]^r[3]^r[1]^g[108]^g[112]^g[118]^g[119];
	g_next[113] = r[55]^r[54]^r[53]^r[52]^r[51]^r[50]^r[49]^r[48]^r[41]^r[39]^r[38]^r[37]^r[36]^r[35]^r[34]^r[32]^r[27]^r[26]^r[23]^r[22]^r[21]^r[20]^r[17]^r[16]^r[13]^r[10]^r[9]^r[7]^r[6]^r[4]^r[3]^r[0]^g[105]^g[109]^g[113]^g[119];
	g_next[114] = r[54]^r[52]^r[50]^r[48]^r[40]^r[39]^r[37]^r[35]^r[33]^r[32]^r[26]^r[22]^r[20]^r[16]^r[12]^r[11]^r[10]^r[8]^r[7]^r[5]^r[4]^r[2]^r[1]^r[0]^g[106]^g[110]^g[114];
	g_next[115] = r[53]^r[52]^r[49]^r[48]^r[39]^r[36]^r[35]^r[32]^r[25]^r[24]^r[23]^r[22]^r[19]^r[18]^r[17]^r[16]^r[11]^r[9]^r[8]^r[6]^r[5]^r[3]^r[2]^r[0]^g[107]^g[111]^g[115];
	g_next[116] = r[52]^r[48]^r[38]^r[37]^r[36]^r[34]^r[33]^r[32]^r[24]^r[22]^r[18]^r[16]^r[10]^r[9]^r[7]^r[6]^r[4]^r[3]^r[1]^r[0]^g[108]^g[112]^g[116];
	g_next[117] = r[51]^r[50]^r[49]^r[48]^r[37]^r[35]^r[34]^r[32]^r[23]^r[22]^r[17]^r[16]^r[9]^r[6]^r[3]^r[0]^g[109]^g[113]^g[117];
	g_next[118] = r[50]^r[48]^r[36]^r[35]^r[33]^r[32]^r[22]^r[16]^r[8]^r[7]^r[6]^r[2]^r[1]^r[0]^g[110]^g[114]^g[118];
	g_next[119] = r[49]^r[48]^r[35]^r[32]^r[21]^r[20]^r[19]^r[18]^r[17]^r[16]^r[7]^r[5]^r[4]^r[3]^r[2]^r[0]^g[111]^g[115]^g[119];
	g_next[120] = r[63]^r[58]^r[56]^r[53]^r[52]^r[50]^r[49]^r[48]^r[44]^r[43]^r[42]^r[41]^r[38]^r[37]^r[35]^r[34]^r[33]^r[30]^r[28]^r[26]^r[25]^r[23]^r[22]^r[21]^r[19]^r[18]^r[16]^r[14]^r[13]^r[12]^r[11]^r[10]^r[7]^r[5]^r[4]^r[3]^r[2]^g[123]^g[125]^g[126]^g[127]^g[129]^g[130];
	g_next[121] = r[58]^r[57]^r[55]^r[52]^r[50]^r[44]^r[43]^r[40]^r[39]^r[38]^r[37]^r[36]^r[34]^r[30]^r[27]^r[25]^r[22]^r[20]^r[16]^r[15]^r[14]^r[11]^r[10]^r[9]^r[8]^r[4]^r[2]^r[1]^g[123]^g[124]^g[125]^g[128]^g[129]^g[131];
	g_next[122] = r[62]^r[57]^r[55]^r[53]^r[51]^r[50]^r[47]^r[43]^r[41]^r[40]^r[39]^r[38]^r[36]^r[34]^r[32]^r[27]^r[24]^r[23]^r[22]^r[17]^r[14]^r[13]^r[8]^r[6]^r[5]^r[4]^r[2]^r[1]^g[124]^g[125]^g[126]^g[129]^g[130]^g[132];
	g_next[123] = r[62]^r[57]^r[54]^r[50]^r[48]^r[47]^r[39]^r[37]^r[36]^r[34]^r[32]^r[29]^r[28]^r[22]^r[20]^r[18]^r[17]^r[13]^r[12]^r[10]^r[8]^r[6]^r[4]^r[2]^r[1]^r[0]^g[125]^g[126]^g[127]^g[130]^g[131]^g[133];
	g_next[124] = r[61]^r[57]^r[52]^r[51]^r[50]^r[46]^r[43]^r[40]^r[36]^r[31]^r[29]^r[24]^r[23]^r[22]^r[19]^r[16]^r[15]^r[14]^r[12]^r[10]^r[9]^r[8]^r[5]^r[4]^g[126]^g[127]^g[128]^g[131]^g[132]^g[134];
	g_next[125] = r[54]^r[53]^r[52]^r[50]^r[47]^r[42]^r[40]^r[39]^r[37]^r[36]^r[28]^r[27]^r[26]^r[23]^r[22]^r[19]^r[17]^r[13]^r[11]^r[9]^r[4]^g[120]^g[127]^g[128]^g[129]^g[132]^g[133];
	g_next[126] = r[61]^r[60]^r[53]^r[51]^r[50]^r[47]^r[46]^r[45]^r[42]^r[39]^r[38]^r[36]^r[33]^r[31]^r[30]^r[27]^r[23]^r[22]^r[19]^r[18]^r[17]^r[16]^r[15]^r[14]^r[13]^r[12]^r[8]^r[5]^r[4]^r[1]^r[0]^g[120]^g[121]^g[128]^g[129]^g[130]^g[133]^g[134];
	g_next[127] = r[60]^r[56]^r[53]^r[52]^r[50]^r[46]^r[45]^r[42]^r[41]^r[38]^r[36]^r[30]^r[28]^r[27]^r[26]^r[25]^r[23]^r[16]^r[15]^r[14]^r[13]^r[12]^r[11]^r[10]^r[9]^r[7]^r[4]^g[121]^g[122]^g[129]^g[130]^g[131]^g[134];
	g_next[128] = r[60]^r[59]^r[53]^r[51]^r[50]^r[45]^r[44]^r[39]^r[37]^r[36]^r[32]^r[30]^r[29]^r[27]^r[25]^r[17]^r[15]^r[14]^r[13]^r[11]^r[10]^r[8]^r[7]^r[4]^r[0]^g[120]^g[122]^g[123]^g[130]^g[131]^g[132];
	g_next[129] = r[60]^r[55]^r[51]^r[50]^r[46]^r[40]^r[38]^r[32]^r[30]^r[27]^r[25]^r[24]^r[21]^r[18]^r[17]^r[16]^r[10]^r[9]^r[8]^r[7]^r[6]^r[4]^r[0]^g[120]^g[121]^g[123]^g[124]^g[131]^g[132]^g[133];
	g_next[130] = r[58]^r[55]^r[51]^r[50]^r[45]^r[43]^r[41]^r[40]^r[38]^r[37]^r[36]^r[31]^r[28]^r[27]^r[25]^r[22]^r[16]^r[15]^r[11]^r[8]^r[7]^g[120]^g[121]^g[122]^g[124]^g[125]^g[132]^g[133]^g[134];
	g_next[131] = r[58]^r[54]^r[52]^r[45]^r[44]^r[43]^r[39]^r[38]^r[37]^r[36]^r[35]^r[28]^r[23]^r[20]^r[17]^r[15]^r[14]^r[13]^r[12]^r[10]^r[8]^r[5]^g[121]^g[122]^g[123]^g[125]^g[126]^g[133]^g[134];
	g_next[132] = r[59]^r[57]^r[45]^r[44]^r[42]^r[40]^r[36]^r[35]^r[31]^r[30]^r[29]^r[27]^r[23]^r[21]^r[20]^r[17]^r[16]^r[14]^r[10]^r[9]^r[8]^r[5]^r[3]^g[120]^g[122]^g[123]^g[124]^g[126]^g[127]^g[134];
	g_next[133] = r[54]^r[53]^r[51]^r[50]^r[49]^r[43]^r[40]^r[39]^r[38]^r[34]^r[30]^r[26]^r[24]^r[22]^r[21]^r[19]^r[16]^r[15]^r[13]^r[12]^r[11]^r[10]^r[9]^r[6]^r[4]^g[121]^g[123]^g[124]^g[125]^g[127]^g[128];
	g_next[134] = r[58]^r[57]^r[56]^r[53]^r[51]^r[42]^r[41]^r[39]^r[38]^r[37]^r[36]^r[30]^r[29]^r[28]^r[27]^r[26]^r[20]^r[15]^r[14]^r[12]^r[11]^r[8]^r[2]^g[122]^g[124]^g[125]^g[126]^g[128]^g[129];
	g_next[135] = r[63]^r[60]^r[57]^r[54]^r[52]^r[51]^r[48]^r[46]^r[45]^r[41]^r[39]^r[38]^r[33]^r[32]^r[30]^r[29]^r[28]^r[27]^r[20]^r[19]^r[15]^r[13]^r[6]^r[3]^r[1]^r[0]^g[138]^g[141]^g[142]^g[145]^g[146]^g[149];
	g_next[136] = r[60]^r[59]^r[52]^r[46]^r[45]^r[44]^r[43]^r[39]^r[37]^r[32]^r[31]^r[29]^r[28]^r[26]^r[23]^r[20]^r[19]^r[18]^r[16]^r[15]^r[7]^r[6]^r[2]^r[1]^r[0]^g[135]^g[138]^g[139]^g[141]^g[143]^g[145]^g[147]^g[149];
	g_next[137] = r[59]^r[57]^r[55]^r[48]^r[45]^r[44]^r[43]^r[42]^r[41]^r[39]^r[37]^r[34]^r[31]^r[27]^r[26]^r[25]^r[22]^r[20]^r[19]^r[18]^r[14]^r[12]^r[11]^r[10]^r[7]^r[4]^r[0]^g[136]^g[139]^g[140]^g[142]^g[144]^g[146]^g[148];
	g_next[138] = r[54]^r[53]^r[52]^r[51]^r[48]^r[45]^r[44]^r[41]^r[40]^r[39]^r[37]^r[36]^r[34]^r[31]^r[30]^r[25]^r[22]^r[21]^r[18]^r[17]^r[16]^r[15]^r[12]^r[10]^r[9]^r[6]^r[4]^r[2]^r[1]^r[0]^g[137]^g[140]^g[141]^g[143]^g[145]^g[147]^g[149];
	g_next[139] = r[62]^r[55]^r[53]^r[47]^r[45]^r[42]^r[41]^r[39]^r[37]^r[34]^r[33]^r[32]^r[31]^r[28]^r[27]^r[26]^r[23]^r[19]^r[18]^r[17]^r[16]^r[14]^r[11]^r[10]^r[9]^r[6]^r[5]^r[2]^r[1]^g[135]^g[138]^g[141]^g[142]^g[144]^g[146]^g[148];
	g_next[140] = r[62]^r[59]^r[58]^r[52]^r[51]^r[48]^r[47]^r[43]^r[42]^r[40]^r[39]^r[34]^r[32]^r[31]^r[30]^r[26]^r[25]^r[22]^r[21]^r[20]^r[19]^r[18]^r[17]^r[16]^r[14]^r[13]^r[10]^r[6]^r[3]^r[2]^r[1]^r[0]^g[135]^g[136]^g[139]^g[142]^g[143]^g[145]^g[147]^g[149];
	g_next[141] = r[59]^r[56]^r[54]^r[51]^r[47]^r[45]^r[41]^r[40]^r[33]^r[31]^r[28]^r[27]^r[26]^r[24]^r[22]^r[21]^r[15]^r[14]^r[13]^r[11]^r[10]^r[9]^r[5]^r[3]^r[1]^r[0]^g[136]^g[137]^g[140]^g[143]^g[144]^g[146]^g[148];
	g_next[142] = r[58]^r[56]^r[54]^r[53]^r[52]^r[51]^r[50]^r[42]^r[41]^r[39]^r[35]^r[29]^r[26]^r[25]^r[20]^r[19]^r[18]^r[16]^r[15]^r[14]^r[13]^r[10]^r[8]^r[6]^r[5]^r[1]^r[0]^g[137]^g[138]^g[141]^g[144]^g[145]^g[147]^g[149];
	g_next[143] = r[61]^r[54]^r[53]^r[51]^r[50]^r[47]^r[46]^r[43]^r[41]^r[39]^r[35]^r[32]^r[31]^r[29]^r[27]^r[26]^r[25]^r[24]^r[22]^r[21]^r[20]^r[18]^r[14]^r[13]^r[11]^r[10]^r[4]^r[3]^g[135]^g[138]^g[139]^g[142]^g[145]^g[146]^g[148];
	g_next[144] = r[58]^r[57]^r[54]^r[52]^r[51]^r[50]^r[47]^r[44]^r[42]^r[40]^r[39]^r[36]^r[32]^r[29]^r[27]^r[26]^r[24]^r[22]^r[21]^r[20]^r[19]^r[12]^r[10]^r[8]^r[4]^r[2]^g[135]^g[136]^g[139]^g[140]^g[143]^g[146]^g[147]^g[149];
	g_next[145] = r[61]^r[57]^r[55]^r[53]^r[51]^r[47]^r[44]^r[42]^r[41]^r[40]^r[38]^r[33]^r[32]^r[31]^r[29]^r[27]^r[26]^r[24]^r[23]^r[19]^r[18]^r[17]^r[16]^r[15]^r[14]^r[10]^r[8]^r[5]^r[4]^r[1]^g[136]^g[137]^g[140]^g[141]^g[144]^g[147]^g[148];
	g_next[146] = r[58]^r[57]^r[52]^r[51]^r[49]^r[46]^r[44]^r[41]^r[39]^r[38]^r[34]^r[32]^r[30]^r[28]^r[27]^r[26]^r[24]^r[23]^r[21]^r[20]^r[19]^r[18]^r[17]^r[15]^r[10]^r[8]^r[7]^r[5]^r[2]^g[137]^g[138]^g[141]^g[142]^g[145]^g[148]^g[149];
	g_next[147] = r[60]^r[57]^r[55]^r[51]^r[46]^r[45]^r[42]^r[41]^r[31]^r[30]^r[26]^r[23]^r[21]^r[20]^r[18]^r[15]^r[14]^r[10]^r[7]^r[5]^r[4]^r[3]^r[2]^r[0]^g[135]^g[138]^g[139]^g[142]^g[143]^g[146]^g[149];
	g_next[148] = r[60]^r[57]^r[56]^r[52]^r[51]^r[45]^r[43]^r[42]^r[41]^r[40]^r[39]^r[35]^r[34]^r[30]^r[24]^r[18]^r[17]^r[13]^r[12]^r[11]^r[10]^r[7]^r[2]^r[1]^g[136]^g[139]^g[140]^g[143]^g[144]^g[147];
	g_next[149] = r[60]^r[57]^r[54]^r[53]^r[52]^r[51]^r[49]^r[40]^r[38]^r[37]^r[35]^r[32]^r[30]^r[22]^r[21]^r[20]^r[19]^r[17]^r[16]^r[15]^r[14]^r[13]^r[11]^r[4]^r[1]^r[0]^g[137]^g[140]^g[141]^g[144]^g[145]^g[148];
	g_next[150] = r[63]^r[58]^r[53]^r[52]^r[48]^r[46]^r[43]^r[41]^r[38]^r[36]^r[33]^r[32]^r[30]^r[29]^r[28]^r[26]^r[23]^r[20]^r[19]^r[13]^r[10]^r[9]^r[8]^r[6]^r[3]^r[1]^r[0]^g[151]^g[153]^g[154]^g[158]^g[159]^g[163]^g[164];
	g_next[151] = r[58]^r[43]^r[41]^r[38]^r[36]^r[32]^r[30]^r[26]^r[24]^r[23]^r[22]^r[20]^r[19]^r[18]^r[16]^r[11]^r[10]^r[8]^r[7]^r[6]^r[4]^r[3]^g[150]^g[151]^g[152]^g[153]^g[155]^g[158]^g[160]^g[163];
	g_next[152] = r[58]^r[54]^r[53]^r[44]^r[43]^r[42]^r[41]^r[34]^r[30]^r[28]^r[20]^r[18]^r[13]^r[11]^r[10]^r[9]^r[7]^r[6]^r[4]^r[3]^r[1]^g[150]^g[151]^g[152]^g[153]^g[154]^g[156]^g[159]^g[161]^g[164];
	g_next[153] = r[60]^r[58]^r[55]^r[54]^r[50]^r[48]^r[45]^r[41]^r[40]^r[36]^r[35]^r[34]^r[31]^r[28]^r[26]^r[25]^r[24]^r[23]^r[21]^r[20]^r[19]^r[18]^r[16]^r[15]^r[12]^r[7]^r[6]^r[5]^r[4]^r[2]^g[151]^g[152]^g[153]^g[154]^g[155]^g[157]^g[160]^g[162];
	g_next[154] = r[58]^r[55]^r[53]^r[50]^r[48]^r[44]^r[43]^r[42]^r[41]^r[35]^r[34]^r[31]^r[28]^r[26]^r[24]^r[15]^r[10]^r[7]^r[4]^r[2]^g[152]^g[153]^g[154]^g[155]^g[156]^g[158]^g[161]^g[163];
	g_next[155] = r[58]^r[56]^r[55]^r[46]^r[44]^r[43]^r[41]^r[40]^r[34]^r[32]^r[28]^r[25]^r[23]^r[22]^r[21]^r[20]^r[19]^r[16]^r[15]^r[8]^r[7]^r[6]^r[4]^r[0]^g[153]^g[154]^g[155]^g[156]^g[157]^g[159]^g[162]^g[164];
	g_next[156] = r[62]^r[58]^r[57]^r[55]^r[54]^r[53]^r[52]^r[50]^r[47]^r[46]^r[45]^r[43]^r[41]^r[38]^r[37]^r[34]^r[33]^r[32]^r[30]^r[27]^r[26]^r[25]^r[23]^r[21]^r[20]^r[17]^r[15]^r[14]^r[12]^r[10]^r[9]^r[6]^r[5]^g[150]^g[154]^g[155]^g[156]^g[157]^g[158]^g[160]^g[163];
	g_next[157] = r[62]^r[60]^r[58]^r[56]^r[54]^r[50]^r[48]^r[47]^r[46]^r[44]^r[42]^r[41]^r[40]^r[38]^r[36]^r[35]^r[34]^r[31]^r[28]^r[27]^r[26]^r[24]^r[22]^r[19]^r[16]^r[15]^r[14]^r[8]^r[6]^r[5]^r[4]^r[2]^g[150]^g[151]^g[155]^g[156]^g[157]^g[158]^g[159]^g[161]^g[164];
	g_next[158] = r[53]^r[52]^r[43]^r[41]^r[37]^r[35]^r[33]^r[31]^r[27]^r[25]^r[23]^r[22]^r[21]^r[18]^r[15]^r[12]^r[8]^r[7]^r[0]^g[151]^g[152]^g[156]^g[157]^g[158]^g[159]^g[160]^g[162];
	g_next[159] = r[59]^r[54]^r[52]^r[49]^r[47]^r[44]^r[43]^r[42]^r[41]^r[39]^r[35]^r[34]^r[30]^r[29]^r[25]^r[24]^r[23]^r[22]^r[20]^r[18]^r[15]^r[14]^r[12]^r[11]^r[10]^r[9]^r[8]^r[4]^r[2]^r[1]^r[0]^g[152]^g[153]^g[157]^g[158]^g[159]^g[160]^g[161]^g[163];
	g_next[160] = r[59]^r[53]^r[52]^r[44]^r[43]^r[42]^r[41]^r[39]^r[35]^r[24]^r[22]^r[20]^r[19]^r[18]^r[17]^r[15]^r[11]^r[9]^r[5]^r[4]^g[153]^g[154]^g[158]^g[159]^g[160]^g[161]^g[162]^g[164];
	g_next[161] = r[55]^r[52]^r[49]^r[47]^r[45]^r[41]^r[39]^r[34]^r[31]^r[30]^r[25]^r[24]^r[23]^r[22]^r[21]^r[20]^r[19]^r[18]^r[15]^r[9]^r[7]^r[5]^r[1]^g[150]^g[154]^g[155]^g[159]^g[160]^g[161]^g[162]^g[163];
	g_next[162] = r[61]^r[56]^r[55]^r[53]^r[52]^r[51]^r[49]^r[46]^r[44]^r[43]^r[39]^r[37]^r[36]^r[32]^r[29]^r[27]^r[26]^r[25]^r[21]^r[18]^r[16]^r[15]^r[13]^r[11]^r[9]^r[8]^r[7]^r[6]^r[4]^r[3]^g[150]^g[151]^g[155]^g[156]^g[160]^g[161]^g[162]^g[163]^g[164];
	g_next[163] = r[59]^r[56]^r[55]^r[54]^r[52]^r[51]^r[47]^r[44]^r[43]^r[42]^r[41]^r[39]^r[36]^r[35]^r[34]^r[32]^r[31]^r[30]^r[29]^r[27]^r[24]^r[23]^r[22]^r[21]^r[20]^r[19]^r[18]^r[16]^r[15]^r[11]^r[9]^r[8]^r[7]^r[3]^r[1]^g[151]^g[152]^g[156]^g[157]^g[161]^g[162]^g[163]^g[164];
	g_next[164] = r[61]^r[59]^r[57]^r[55]^r[53]^r[52]^r[51]^r[49]^r[47]^r[46]^r[45]^r[43]^r[42]^r[41]^r[39]^r[37]^r[36]^r[35]^r[33]^r[32]^r[27]^r[25]^r[24]^r[23]^r[22]^r[20]^r[18]^r[17]^r[15]^r[13]^r[11]^r[6]^r[5]^r[4]^r[3]^r[1]^g[150]^g[152]^g[153]^g[157]^g[158]^g[162]^g[163]^g[164];
	g_next[165] = r[63]^r[58]^r[53]^r[52]^r[48]^r[43]^r[41]^r[38]^r[36]^r[33]^r[32]^r[30]^r[28]^r[23]^r[20]^r[19]^r[18]^r[14]^r[13]^r[12]^r[10]^r[9]^r[4]^r[3]^r[1]^r[0]^g[168]^g[170]^g[172]^g[174]^g[179];
	g_next[166] = r[61]^r[55]^r[54]^r[52]^r[50]^r[47]^r[46]^r[43]^r[38]^r[31]^r[27]^r[26]^r[23]^r[22]^r[20]^r[18]^r[16]^r[12]^r[11]^r[10]^r[9]^r[7]^r[5]^r[4]^r[3]^r[1]^r[0]^g[165]^g[168]^g[169]^g[170]^g[171]^g[172]^g[173]^g[174]^g[175]^g[179];
	g_next[167] = r[61]^r[59]^r[55]^r[48]^r[46]^r[45]^r[43]^r[41]^r[37]^r[34]^r[29]^r[28]^r[27]^r[16]^r[14]^r[13]^r[12]^r[11]^r[9]^r[8]^r[7]^r[5]^r[3]^r[2]^r[1]^g[166]^g[169]^g[170]^g[171]^g[172]^g[173]^g[174]^g[175]^g[176];
	g_next[168] = r[61]^r[58]^r[57]^r[54]^r[50]^r[48]^r[45]^r[44]^r[43]^r[42]^r[39]^r[34]^r[33]^r[31]^r[30]^r[29]^r[28]^r[27]^r[26]^r[25]^r[24]^r[23]^r[20]^r[16]^r[14]^r[13]^r[9]^r[6]^r[2]^g[167]^g[170]^g[171]^g[172]^g[173]^g[174]^g[175]^g[176]^g[177];
	g_next[169] = r[61]^r[59]^r[57]^r[56]^r[55]^r[50]^r[48]^r[47]^r[46]^r[45]^r[43]^r[40]^r[39]^r[31]^r[26]^r[25]^r[24]^r[19]^r[14]^r[13]^r[11]^r[10]^r[9]^r[6]^r[5]^r[4]^r[2]^r[0]^g[168]^g[171]^g[172]^g[173]^g[174]^g[175]^g[176]^g[177]^g[178];
	g_next[170] = r[56]^r[54]^r[53]^r[50]^r[48]^r[46]^r[44]^r[43]^r[42]^r[40]^r[39]^r[38]^r[36]^r[35]^r[31]^r[29]^r[28]^r[25]^r[24]^r[20]^r[17]^r[16]^r[14]^r[12]^r[11]^r[9]^r[6]^r[3]^r[0]^g[169]^g[172]^g[173]^g[174]^g[175]^g[176]^g[177]^g[178]^g[179];
	g_next[171] = r[59]^r[56]^r[51]^r[48]^r[45]^r[44]^r[43]^r[39]^r[37]^r[36]^r[35]^r[34]^r[33]^r[31]^r[29]^r[28]^r[27]^r[26]^r[23]^r[22]^r[21]^r[17]^r[15]^r[14]^r[11]^r[9]^r[8]^r[6]^r[5]^r[4]^r[2]^r[0]^g[165]^g[170]^g[173]^g[174]^g[175]^g[176]^g[177]^g[178]^g[179];
	g_next[172] = r[56]^r[54]^r[53]^r[51]^r[49]^r[48]^r[45]^r[43]^r[42]^r[36]^r[35]^r[28]^r[27]^r[26]^r[24]^r[23]^r[22]^r[20]^r[19]^r[17]^r[13]^r[10]^r[9]^r[8]^r[6]^r[1]^r[0]^g[166]^g[171]^g[174]^g[175]^g[176]^g[177]^g[178]^g[179];
	g_next[173] = r[62]^r[59]^r[55]^r[53]^r[47]^r[45]^r[43]^r[37]^r[36]^r[35]^r[34]^r[33]^r[32]^r[31]^r[29]^r[26]^r[24]^r[22]^r[19]^r[15]^r[14]^r[13]^r[12]^r[10]^r[9]^r[1]^g[165]^g[167]^g[172]^g[175]^g[176]^g[177]^g[178]^g[179];
	g_next[174] = r[62]^r[60]^r[54]^r[53]^r[51]^r[48]^r[47]^r[46]^r[45]^r[44]^r[43]^r[38]^r[36]^r[30]^r[29]^r[27]^r[26]^r[24]^r[23]^r[22]^r[20]^r[19]^r[15]^r[14]^r[12]^r[4]^r[3]^r[2]^r[1]^r[0]^g[166]^g[168]^g[173]^g[176]^g[177]^g[178]^g[179];
	g_next[175] = r[58]^r[53]^r[51]^r[49]^r[47]^r[46]^r[44]^r[40]^r[37]^r[36]^r[33]^r[30]^r[28]^r[27]^r[25]^r[22]^r[21]^r[19]^r[17]^r[13]^r[12]^r[9]^r[7]^r[3]^r[1]^g[165]^g[167]^g[169]^g[174]^g[177]^g[178]^g[179];
	g_next[176] = r[58]^r[57]^r[56]^r[54]^r[53]^r[49]^r[45]^r[43]^r[41]^r[40]^r[38]^r[36]^r[32]^r[30]^r[29]^r[25]^r[24]^r[23]^r[22]^r[19]^r[11]^r[10]^r[7]^r[6]^r[5]^r[4]^r[2]^r[0]^g[166]^g[168]^g[170]^g[175]^g[178]^g[179];
	g_next[177] = r[58]^r[57]^r[55]^r[54]^r[53]^r[46]^r[45]^r[43]^r[41]^r[39]^r[33]^r[32]^r[29]^r[28]^r[27]^r[26]^r[22]^r[19]^r[18]^r[15]^r[10]^r[9]^r[4]^r[3]^g[165]^g[167]^g[169]^g[171]^g[176]^g[179];
	g_next[178] = r[60]^r[58]^r[56]^r[54]^r[53]^r[52]^r[46]^r[44]^r[43]^r[41]^r[37]^r[35]^r[34]^r[28]^r[27]^r[25]^r[19]^r[18]^r[16]^r[15]^r[12]^r[11]^r[9]^r[4]^r[3]^r[2]^r[1]^g[166]^g[168]^g[170]^g[172]^g[177];
	g_next[179] = r[58]^r[53]^r[52]^r[50]^r[49]^r[45]^r[44]^r[41]^r[39]^r[37]^r[36]^r[33]^r[32]^r[26]^r[25]^r[24]^r[23]^r[22]^r[21]^r[20]^r[19]^r[15]^r[14]^r[11]^r[7]^r[4]^r[3]^r[2]^r[1]^g[167]^g[169]^g[171]^g[173]^g[178];
	g_next[180] = r[63]^r[60]^r[57]^r[51]^r[48]^r[46]^r[44]^r[42]^r[40]^r[39]^r[38]^r[33]^r[30]^r[29]^r[28]^r[25]^r[24]^r[21]^r[17]^r[16]^r[15]^r[13]^r[4]^r[3]^r[2]^g[182]^g[183]^g[184]^g[185]^g[187]^g[188]^g[189]^g[190]^g[191]^g[194];
	g_next[181] = r[60]^r[59]^r[51]^r[46]^r[45]^r[42]^r[41]^r[40]^r[38]^r[36]^r[35]^r[33]^r[32]^r[31]^r[28]^r[26]^r[24]^r[23]^r[18]^r[16]^r[15]^r[12]^r[7]^r[6]^r[5]^r[4]^r[3]^r[2]^g[180]^g[182]^g[186]^g[187]^g[192]^g[194];
	g_next[182] = r[59]^r[57]^r[55]^r[54]^r[51]^r[50]^r[46]^r[45]^r[41]^r[39]^r[36]^r[35]^r[33]^r[32]^r[31]^r[29]^r[27]^r[26]^r[23]^r[22]^r[21]^r[19]^r[18]^r[17]^r[16]^r[15]^r[14]^r[13]^r[10]^r[9]^r[5]^r[1]^r[0]^g[181]^g[183]^g[187]^g[188]^g[193];
	g_next[183] = r[56]^r[54]^r[50]^r[48]^r[47]^r[45]^r[41]^r[38]^r[35]^r[30]^r[29]^r[27]^r[23]^r[22]^r[18]^r[17]^r[16]^r[13]^r[12]^r[7]^g[182]^g[184]^g[188]^g[189]^g[194];
	g_next[184] = r[60]^r[55]^r[54]^r[51]^r[41]^r[39]^r[37]^r[35]^r[32]^r[30]^r[28]^r[26]^r[24]^r[23]^r[19]^r[18]^r[17]^r[16]^r[15]^r[14]^r[13]^r[9]^r[8]^r[4]^r[3]^r[1]^g[180]^g[183]^g[185]^g[189]^g[190];
	g_next[185] = r[61]^r[60]^r[58]^r[55]^r[54]^r[52]^r[51]^r[49]^r[47]^r[45]^r[43]^r[40]^r[37]^r[35]^r[34]^r[32]^r[31]^r[29]^r[28]^r[25]^r[24]^r[23]^r[22]^r[19]^r[15]^r[13]^r[9]^r[8]^r[5]^r[1]^g[180]^g[181]^g[184]^g[186]^g[190]^g[191];
	g_next[186] = r[61]^r[55]^r[54]^r[52]^r[51]^r[47]^r[46]^r[43]^r[42]^r[36]^r[35]^r[34]^r[33]^r[30]^r[29]^r[28]^r[27]^r[26]^r[25]^r[23]^r[18]^r[15]^r[14]^r[9]^r[7]^r[6]^r[5]^r[1]^r[0]^g[180]^g[181]^g[182]^g[185]^g[187]^g[191]^g[192];
	g_next[187] = r[61]^r[56]^r[54]^r[49]^r[46]^r[45]^r[43]^r[42]^r[36]^r[35]^r[33]^r[31]^r[30]^r[29]^r[27]^r[25]^r[20]^r[18]^r[17]^r[16]^r[14]^r[13]^r[11]^r[10]^r[9]^r[8]^r[6]^r[5]^r[2]^g[180]^g[181]^g[182]^g[183]^g[186]^g[188]^g[192]^g[193];
	g_next[188] = r[61]^r[57]^r[54]^r[52]^r[49]^r[48]^r[47]^r[43]^r[39]^r[35]^r[34]^r[33]^r[31]^r[29]^r[27]^r[26]^r[25]^r[24]^r[19]^r[17]^r[15]^r[13]^r[9]^r[8]^r[7]^r[6]^r[5]^r[1]^r[0]^g[180]^g[181]^g[182]^g[183]^g[184]^g[187]^g[189]^g[193]^g[194];
	g_next[189] = r[55]^r[54]^r[52]^r[49]^r[46]^r[45]^r[43]^r[40]^r[38]^r[35]^r[30]^r[24]^r[19]^r[15]^r[13]^r[11]^r[8]^r[6]^r[4]^r[0]^g[181]^g[182]^g[183]^g[184]^g[185]^g[188]^g[190]^g[194];
	g_next[190] = r[62]^r[59]^r[57]^r[56]^r[55]^r[54]^r[53]^r[50]^r[49]^r[47]^r[46]^r[44]^r[43]^r[41]^r[39]^r[38]^r[36]^r[34]^r[32]^r[31]^r[30]^r[27]^r[23]^r[20]^r[19]^r[17]^r[16]^r[15]^r[14]^r[13]^r[10]^r[8]^r[7]^r[5]^r[2]^r[1]^g[180]^g[182]^g[183]^g[184]^g[185]^g[186]^g[189]^g[191];
	g_next[191] = r[62]^r[56]^r[54]^r[53]^r[49]^r[48]^r[47]^r[46]^r[45]^r[44]^r[40]^r[38]^r[37]^r[36]^r[34]^r[31]^r[29]^r[28]^r[27]^r[26]^r[16]^r[13]^r[11]^r[10]^r[7]^r[4]^r[2]^r[1]^g[180]^g[181]^g[183]^g[184]^g[185]^g[186]^g[187]^g[190]^g[192];
	g_next[192] = r[59]^r[56]^r[54]^r[53]^r[49]^r[41]^r[39]^r[38]^r[37]^r[28]^r[27]^r[26]^r[23]^r[21]^r[20]^r[18]^r[16]^r[13]^r[12]^r[11]^r[9]^r[8]^r[6]^r[5]^r[3]^r[2]^r[1]^r[0]^g[180]^g[181]^g[182]^g[184]^g[185]^g[186]^g[187]^g[188]^g[191]^g[193];
	g_next[193] = r[58]^r[56]^r[55]^r[54]^r[50]^r[47]^r[46]^r[45]^r[38]^r[37]^r[35]^r[32]^r[31]^r[30]^r[29]^r[25]^r[20]^r[18]^r[14]^r[13]^r[11]^r[9]^r[8]^r[6]^r[4]^r[0]^g[180]^g[181]^g[182]^g[183]^g[185]^g[186]^g[187]^g[188]^g[189]^g[192]^g[194];
	g_next[194] = r[59]^r[55]^r[54]^r[50]^r[49]^r[47]^r[46]^r[44]^r[38]^r[37]^r[36]^r[31]^r[28]^r[27]^r[26]^r[25]^r[23]^r[21]^r[18]^r[14]^r[13]^r[11]^r[8]^r[7]^r[6]^r[3]^r[2]^r[0]^g[181]^g[182]^g[183]^g[184]^g[186]^g[187]^g[188]^g[189]^g[190]^g[193];
	g_next[195] = r[63]^r[58]^r[53]^r[52]^r[50]^r[48]^r[43]^r[42]^r[41]^r[40]^r[37]^r[36]^r[33]^r[32]^r[30]^r[26]^r[24]^r[23]^r[22]^r[21]^r[20]^r[19]^r[18]^r[17]^r[14]^r[12]^r[11]^r[10]^r[9]^r[6]^r[4]^r[3]^r[1]^r[0]^g[196]^g[197]^g[198]^g[199]^g[200]^g[201]^g[203]^g[205]^g[209];
	g_next[196] = r[58]^r[55]^r[53]^r[52]^r[51]^r[50]^r[47]^r[46]^r[42]^r[38]^r[37]^r[36]^r[33]^r[31]^r[30]^r[29]^r[28]^r[27]^r[26]^r[24]^r[23]^r[20]^r[17]^r[11]^r[10]^r[7]^r[6]^r[4]^r[3]^r[2]^r[1]^g[195]^g[196]^g[202]^g[203]^g[204]^g[205]^g[206]^g[209];
	g_next[197] = r[56]^r[55]^r[52]^r[51]^r[48]^r[46]^r[43]^r[41]^r[39]^r[38]^r[33]^r[32]^r[30]^r[28]^r[27]^r[26]^r[24]^r[23]^r[21]^r[17]^r[13]^r[12]^r[9]^r[7]^r[2]^r[1]^r[0]^g[196]^g[197]^g[203]^g[204]^g[205]^g[206]^g[207];
	g_next[198] = r[59]^r[56]^r[55]^r[54]^r[53]^r[52]^r[49]^r[48]^r[46]^r[44]^r[42]^r[39]^r[37]^r[34]^r[32]^r[31]^r[30]^r[28]^r[26]^r[25]^r[22]^r[20]^r[19]^r[18]^r[17]^r[15]^r[11]^r[10]^r[9]^r[5]^r[4]^r[0]^g[197]^g[198]^g[204]^g[205]^g[206]^g[207]^g[208];
	g_next[199] = r[59]^r[55]^r[54]^r[53]^r[47]^r[46]^r[41]^r[37]^r[34]^r[33]^r[31]^r[29]^r[26]^r[25]^r[23]^r[18]^r[17]^r[13]^r[11]^r[9]^r[8]^r[5]^r[4]^r[3]^r[1]^g[198]^g[199]^g[205]^g[206]^g[207]^g[208]^g[209];
	g_next[200] = r[59]^r[57]^r[55]^r[54]^r[48]^r[47]^r[46]^r[40]^r[37]^r[33]^r[32]^r[30]^r[29]^r[27]^r[26]^r[24]^r[20]^r[19]^r[17]^r[15]^r[14]^r[13]^r[11]^r[9]^r[8]^r[5]^r[4]^r[3]^r[2]^r[1]^r[0]^g[195]^g[199]^g[200]^g[206]^g[207]^g[208]^g[209];
	g_next[201] = r[60]^r[59]^r[57]^r[56]^r[50]^r[49]^r[46]^r[45]^r[43]^r[41]^r[40]^r[38]^r[37]^r[35]^r[34]^r[32]^r[27]^r[25]^r[21]^r[20]^r[19]^r[17]^r[16]^r[13]^r[12]^r[10]^r[9]^r[8]^r[6]^r[4]^r[3]^g[196]^g[200]^g[201]^g[207]^g[208]^g[209];
	g_next[202] = r[60]^r[59]^r[57]^r[56]^r[46]^r[42]^r[40]^r[38]^r[37]^r[35]^r[34]^r[33]^r[29]^r[20]^r[18]^r[17]^r[15]^r[13]^r[12]^r[11]^r[10]^r[8]^r[6]^r[3]^r[1]^r[0]^g[195]^g[197]^g[201]^g[202]^g[208]^g[209];
	g_next[203] = r[59]^r[58]^r[57]^r[55]^r[50]^r[48]^r[47]^r[46]^r[45]^r[43]^r[40]^r[37]^r[35]^r[33]^r[32]^r[31]^r[30]^r[28]^r[19]^r[18]^r[17]^r[15]^r[14]^r[13]^r[8]^r[5]^r[2]^r[1]^r[0]^g[196]^g[198]^g[202]^g[203]^g[209];
	g_next[204] = r[61]^r[59]^r[58]^r[56]^r[51]^r[50]^r[47]^r[44]^r[41]^r[40]^r[39]^r[37]^r[36]^r[34]^r[29]^r[28]^r[26]^r[22]^r[21]^r[15]^r[14]^r[12]^r[9]^r[8]^r[7]^r[6]^r[5]^r[4]^r[3]^r[1]^r[0]^g[195]^g[197]^g[199]^g[203]^g[204];
	g_next[205] = r[61]^r[60]^r[59]^r[55]^r[50]^r[48]^r[46]^r[45]^r[41]^r[40]^r[39]^r[38]^r[37]^r[36]^r[34]^r[33]^r[32]^r[31]^r[28]^r[21]^r[17]^r[16]^r[15]^r[12]^r[11]^r[9]^r[8]^r[7]^r[5]^r[4]^g[195]^g[196]^g[198]^g[200]^g[204]^g[205];
	g_next[206] = r[61]^r[60]^r[50]^r[49]^r[48]^r[46]^r[40]^r[39]^r[38]^r[37]^r[33]^r[32]^r[31]^r[28]^r[26]^r[22]^r[21]^r[20]^r[19]^r[18]^r[16]^r[12]^r[8]^r[7]^r[5]^r[4]^r[2]^r[0]^g[195]^g[196]^g[197]^g[199]^g[201]^g[205]^g[206];
	g_next[207] = r[62]^r[61]^r[57]^r[55]^r[52]^r[51]^r[50]^r[46]^r[42]^r[39]^r[36]^r[35]^r[34]^r[33]^r[32]^r[31]^r[30]^r[29]^r[28]^r[27]^r[23]^r[22]^r[21]^r[17]^r[13]^r[12]^r[11]^r[10]^r[6]^r[2]^r[1]^r[0]^g[195]^g[196]^g[197]^g[198]^g[200]^g[202]^g[206]^g[207];
	g_next[208] = r[62]^r[56]^r[51]^r[50]^r[48]^r[47]^r[42]^r[41]^r[35]^r[34]^r[31]^r[29]^r[28]^r[26]^r[21]^r[20]^r[19]^r[17]^r[13]^r[10]^r[9]^r[7]^r[6]^r[4]^r[2]^g[195]^g[196]^g[197]^g[198]^g[199]^g[201]^g[203]^g[207]^g[208];
	g_next[209] = r[57]^r[55]^r[52]^r[49]^r[47]^r[46]^r[42]^r[41]^r[40]^r[38]^r[36]^r[35]^r[31]^r[30]^r[28]^r[20]^r[19]^r[12]^r[11]^r[10]^r[9]^r[8]^r[5]^r[3]^r[2]^g[195]^g[196]^g[197]^g[198]^g[199]^g[200]^g[202]^g[204]^g[208]^g[209];
	g_next[210] = r[63]^r[62]^r[61]^r[59]^r[55]^r[47]^r[46]^r[34]^r[31]^r[30]^r[29]^r[28]^r[22]^r[20]^r[16]^r[14]^r[12]^r[8]^r[5]^r[4]^r[0]^g[210]^g[212]^g[215]^g[218]^g[219]^g[222]^g[223];
	g_next[211] = r[62]^r[60]^r[56]^r[49]^r[48]^r[46]^r[43]^r[41]^r[39]^r[33]^r[32]^r[31]^r[30]^r[20]^r[18]^r[17]^r[16]^r[13]^r[12]^r[8]^r[4]^r[2]^g[211]^g[212]^g[213]^g[215]^g[216]^g[218]^g[220]^g[222]^g[224];
	g_next[212] = r[61]^r[57]^r[50]^r[46]^r[44]^r[43]^r[42]^r[41]^r[40]^r[39]^r[35]^r[34]^r[32]^r[31]^r[29]^r[23]^r[20]^r[19]^r[17]^r[16]^r[15]^r[14]^r[13]^r[12]^r[8]^r[6]^r[4]^r[3]^r[2]^r[1]^r[0]^g[210]^g[212]^g[213]^g[214]^g[216]^g[217]^g[219]^g[221]^g[223];
	g_next[213] = r[60]^r[58]^r[56]^r[51]^r[49]^r[48]^r[47]^r[46]^r[45]^r[44]^r[42]^r[40]^r[39]^r[36]^r[35]^r[31]^r[24]^r[21]^r[15]^r[14]^r[12]^r[9]^r[8]^r[7]^r[5]^r[3]^r[1]^r[0]^g[210]^g[211]^g[213]^g[214]^g[215]^g[217]^g[218]^g[220]^g[222]^g[224];
	g_next[214] = r[59]^r[52]^r[49]^r[48]^r[47]^r[45]^r[44]^r[42]^r[39]^r[37]^r[36]^r[35]^r[34]^r[31]^r[29]^r[25]^r[23]^r[22]^r[20]^r[19]^r[17]^r[14]^r[12]^r[10]^r[9]^r[3]^g[211]^g[212]^g[214]^g[215]^g[216]^g[218]^g[219]^g[221]^g[223];
	g_next[215] = r[58]^r[56]^r[53]^r[51]^r[50]^r[47]^r[44]^r[43]^r[42]^r[39]^r[38]^r[37]^r[32]^r[31]^r[30]^r[26]^r[23]^r[20]^r[18]^r[14]^r[13]^r[12]^r[11]^r[10]^r[9]^r[8]^r[7]^r[5]^r[4]^r[3]^r[1]^r[0]^g[212]^g[213]^g[215]^g[216]^g[217]^g[219]^g[220]^g[222]^g[224];
	g_next[216] = r[57]^r[54]^r[51]^r[49]^r[47]^r[43]^r[42]^r[40]^r[38]^r[37]^r[36]^r[35]^r[34]^r[33]^r[32]^r[29]^r[27]^r[25]^r[24]^r[23]^r[22]^r[21]^r[20]^r[17]^r[15]^r[13]^r[11]^r[8]^r[6]^r[5]^r[4]^r[3]^r[2]^r[1]^g[210]^g[213]^g[214]^g[216]^g[217]^g[218]^g[220]^g[221]^g[223];
	g_next[217] = r[56]^r[55]^r[53]^r[52]^r[51]^r[48]^r[47]^r[42]^r[41]^r[36]^r[35]^r[34]^r[33]^r[32]^r[31]^r[28]^r[25]^r[24]^r[22]^r[21]^r[20]^r[16]^r[13]^r[11]^r[10]^r[8]^r[6]^r[2]^r[1]^g[210]^g[211]^g[214]^g[215]^g[217]^g[218]^g[219]^g[221]^g[222]^g[224];
	g_next[218] = r[56]^r[53]^r[52]^r[51]^r[48]^r[47]^r[40]^r[38]^r[27]^r[26]^r[24]^r[20]^r[15]^r[14]^r[13]^r[12]^r[9]^r[8]^r[7]^r[6]^r[5]^r[4]^r[1]^r[0]^g[211]^g[212]^g[215]^g[216]^g[218]^g[219]^g[220]^g[222]^g[223];
	g_next[219] = r[57]^r[56]^r[55]^r[54]^r[51]^r[49]^r[47]^r[42]^r[39]^r[36]^r[35]^r[34]^r[33]^r[32]^r[31]^r[27]^r[24]^r[22]^r[20]^r[15]^r[14]^r[11]^r[9]^r[7]^r[5]^g[212]^g[213]^g[216]^g[217]^g[219]^g[220]^g[221]^g[223]^g[224];
	g_next[220] = r[58]^r[57]^r[55]^r[53]^r[51]^r[50]^r[47]^r[43]^r[38]^r[37]^r[36]^r[35]^r[34]^r[33]^r[32]^r[28]^r[27]^r[26]^r[25]^r[24]^r[23]^r[21]^r[20]^r[16]^r[14]^r[13]^r[10]^r[9]^r[7]^r[5]^r[4]^r[1]^r[0]^g[210]^g[213]^g[214]^g[217]^g[218]^g[220]^g[221]^g[222]^g[224];
	g_next[221] = r[59]^r[58]^r[57]^r[55]^r[52]^r[49]^r[48]^r[47]^r[44]^r[42]^r[38]^r[37]^r[32]^r[31]^r[29]^r[28]^r[26]^r[25]^r[21]^r[20]^r[17]^r[10]^r[9]^r[8]^r[7]^r[6]^r[2]^r[1]^r[0]^g[211]^g[214]^g[215]^g[218]^g[219]^g[221]^g[222]^g[223];
	g_next[222] = r[60]^r[59]^r[57]^r[56]^r[55]^r[51]^r[49]^r[48]^r[47]^r[45]^r[39]^r[37]^r[36]^r[35]^r[34]^r[30]^r[29]^r[28]^r[25]^r[24]^r[23]^r[22]^r[20]^r[18]^r[16]^r[14]^r[13]^r[11]^r[8]^r[5]^r[4]^r[3]^r[2]^r[0]^g[212]^g[215]^g[216]^g[219]^g[220]^g[222]^g[223]^g[224];
	g_next[223] = r[61]^r[60]^r[59]^r[56]^r[55]^r[50]^r[47]^r[46]^r[44]^r[42]^r[40]^r[36]^r[35]^r[32]^r[30]^r[28]^r[24]^r[23]^r[20]^r[19]^r[15]^r[14]^r[12]^r[10]^r[8]^r[7]^r[5]^r[4]^r[3]^r[2]^r[0]^g[210]^g[213]^g[216]^g[217]^g[220]^g[221]^g[223]^g[224];
	g_next[224] = r[62]^r[61]^r[59]^r[55]^r[49]^r[43]^r[41]^r[39]^r[35]^r[34]^r[33]^r[31]^r[30]^r[28]^r[23]^r[22]^r[21]^r[18]^r[15]^r[14]^r[9]^r[6]^r[2]^r[1]^g[211]^g[214]^g[217]^g[218]^g[221]^g[222]^g[224];
	g_next[225] = r[63]^r[58]^r[56]^r[53]^r[49]^r[44]^r[43]^r[42]^r[40]^r[36]^r[35]^r[30]^r[26]^r[25]^r[24]^r[23]^r[21]^r[20]^r[17]^r[16]^r[12]^r[9]^r[8]^r[7]^r[4]^r[2]^g[228]^g[230]^g[231]^g[232]^g[234]^g[235]^g[236]^g[238]^g[239];
	g_next[226] = r[62]^r[58]^r[56]^r[52]^r[50]^r[48]^r[47]^r[44]^r[42]^r[39]^r[38]^r[37]^r[34]^r[33]^r[32]^r[30]^r[29]^r[26]^r[25]^r[24]^r[23]^r[20]^r[19]^r[18]^r[17]^r[16]^r[14]^r[12]^r[11]^r[10]^r[9]^r[7]^r[4]^r[2]^g[225]^g[228]^g[229]^g[230]^g[233]^g[234]^g[237]^g[238];
	g_next[227] = r[61]^r[56]^r[53]^r[52]^r[49]^r[47]^r[46]^r[41]^r[39]^r[38]^r[36]^r[34]^r[31]^r[29]^r[28]^r[24]^r[23]^r[21]^r[19]^r[17]^r[16]^r[15]^r[13]^r[9]^r[8]^r[7]^r[5]^r[4]^r[3]^r[2]^r[1]^g[225]^g[226]^g[229]^g[230]^g[231]^g[234]^g[235]^g[238]^g[239];
	g_next[228] = r[62]^r[60]^r[57]^r[56]^r[52]^r[50]^r[49]^r[47]^r[46]^r[45]^r[37]^r[36]^r[33]^r[30]^r[29]^r[28]^r[27]^r[25]^r[23]^r[20]^r[19]^r[18]^r[16]^r[15]^r[12]^r[5]^r[3]^r[1]^r[0]^g[226]^g[227]^g[230]^g[231]^g[232]^g[235]^g[236]^g[239];
	g_next[229] = r[59]^r[57]^r[56]^r[48]^r[47]^r[45]^r[44]^r[43]^r[41]^r[38]^r[37]^r[35]^r[33]^r[31]^r[27]^r[26]^r[25]^r[23]^r[16]^r[14]^r[13]^r[10]^r[9]^r[8]^r[6]^r[4]^r[3]^r[2]^r[1]^r[0]^g[225]^g[227]^g[228]^g[231]^g[232]^g[233]^g[236]^g[237];
	g_next[230] = r[60]^r[58]^r[56]^r[52]^r[51]^r[48]^r[47]^r[45]^r[44]^r[43]^r[42]^r[38]^r[36]^r[35]^r[34]^r[33]^r[32]^r[28]^r[27]^r[26]^r[25]^r[24]^r[23]^r[20]^r[18]^r[16]^r[14]^r[13]^r[9]^r[6]^r[5]^r[4]^g[225]^g[226]^g[228]^g[229]^g[232]^g[233]^g[234]^g[237]^g[238];
	g_next[231] = r[61]^r[57]^r[56]^r[50]^r[49]^r[48]^r[47]^r[45]^r[43]^r[42]^r[41]^r[37]^r[36]^r[34]^r[33]^r[31]^r[29]^r[28]^r[25]^r[23]^r[18]^r[14]^r[13]^r[12]^r[11]^r[8]^r[5]^r[3]^r[2]^r[0]^g[225]^g[226]^g[227]^g[229]^g[230]^g[233]^g[234]^g[235]^g[238]^g[239];
	g_next[232] = r[60]^r[58]^r[49]^r[48]^r[43]^r[41]^r[37]^r[35]^r[34]^r[33]^r[28]^r[27]^r[26]^r[25]^r[17]^r[15]^r[11]^r[10]^r[9]^r[8]^r[5]^r[4]^r[3]^r[0]^g[226]^g[227]^g[228]^g[230]^g[231]^g[234]^g[235]^g[236]^g[239];
	g_next[233] = r[55]^r[51]^r[50]^r[48]^r[46]^r[44]^r[43]^r[41]^r[40]^r[37]^r[36]^r[35]^r[31]^r[23]^r[22]^r[19]^r[17]^r[16]^r[15]^r[14]^r[13]^r[12]^r[10]^r[9]^r[7]^r[5]^r[2]^g[225]^g[227]^g[228]^g[229]^g[231]^g[232]^g[235]^g[236]^g[237];
	g_next[234] = r[60]^r[56]^r[55]^r[54]^r[50]^r[48]^r[46]^r[45]^r[44]^r[43]^r[41]^r[39]^r[34]^r[33]^r[32]^r[28]^r[27]^r[24]^r[21]^r[18]^r[17]^r[16]^r[15]^r[14]^r[10]^r[9]^r[8]^r[7]^r[6]^r[2]^g[225]^g[226]^g[228]^g[229]^g[230]^g[232]^g[233]^g[236]^g[237]^g[238];
	g_next[235] = r[57]^r[55]^r[54]^r[53]^r[49]^r[48]^r[45]^r[44]^r[43]^r[38]^r[36]^r[34]^r[31]^r[25]^r[24]^r[23]^r[20]^r[17]^r[15]^r[13]^r[10]^r[6]^r[5]^r[4]^r[3]^r[2]^r[1]^g[225]^g[226]^g[227]^g[229]^g[230]^g[231]^g[233]^g[234]^g[237]^g[238]^g[239];
	g_next[236] = r[56]^r[53]^r[52]^r[50]^r[49]^r[48]^r[45]^r[44]^r[40]^r[39]^r[37]^r[36]^r[34]^r[33]^r[24]^r[23]^r[21]^r[19]^r[18]^r[15]^r[13]^r[11]^r[8]^r[6]^r[5]^r[3]^r[2]^r[0]^g[226]^g[227]^g[228]^g[230]^g[231]^g[232]^g[234]^g[235]^g[238]^g[239];
	g_next[237] = r[59]^r[54]^r[53]^r[52]^r[51]^r[48]^r[45]^r[42]^r[40]^r[39]^r[36]^r[35]^r[31]^r[27]^r[26]^r[22]^r[18]^r[16]^r[15]^r[13]^r[12]^r[10]^r[9]^r[8]^r[6]^r[4]^r[2]^g[225]^g[227]^g[228]^g[229]^g[231]^g[232]^g[233]^g[235]^g[236]^g[239];
	g_next[238] = r[58]^r[56]^r[54]^r[51]^r[50]^r[48]^r[43]^r[42]^r[41]^r[39]^r[38]^r[37]^r[34]^r[33]^r[26]^r[25]^r[24]^r[23]^r[22]^r[21]^r[19]^r[17]^r[16]^r[15]^r[11]^r[8]^r[7]^r[4]^r[2]^r[0]^g[226]^g[228]^g[229]^g[230]^g[232]^g[233]^g[234]^g[236]^g[237];
	g_next[239] = r[57]^r[53]^r[52]^r[51]^r[50]^r[48]^r[44]^r[43]^r[42]^r[41]^r[40]^r[39]^r[37]^r[35]^r[25]^r[24]^r[21]^r[17]^r[16]^r[15]^r[12]^r[6]^r[5]^r[4]^r[3]^r[2]^g[227]^g[229]^g[230]^g[231]^g[233]^g[234]^g[235]^g[237]^g[238];
	g_next[240] = r[63]^r[60]^r[58]^r[57]^r[56]^r[54]^r[53]^r[51]^r[50]^r[49]^r[48]^r[46]^r[45]^r[44]^r[43]^r[42]^r[40]^r[39]^r[38]^r[37]^r[36]^r[35]^r[34]^r[33]^r[32]^r[29]^r[28]^r[27]^r[25]^r[24]^r[23]^r[22]^r[21]^r[17]^r[15]^r[13]^r[11]^r[10]^r[9]^r[7]^r[5]^r[4]^r[3]^r[2]^r[1]^g[245]^g[247]^g[249]^g[253]^g[254];
	g_next[241] = r[60]^r[58]^r[54]^r[53]^r[51]^r[50]^r[49]^r[48]^r[46]^r[43]^r[42]^r[36]^r[35]^r[34]^r[32]^r[29]^r[28]^r[24]^r[20]^r[15]^r[14]^r[12]^r[11]^r[10]^r[9]^r[8]^r[6]^r[4]^r[3]^r[2]^g[240]^g[245]^g[246]^g[247]^g[248]^g[249]^g[250]^g[253];
	g_next[242] = r[58]^r[57]^r[54]^r[51]^r[50]^r[49]^r[48]^r[45]^r[42]^r[39]^r[37]^r[36]^r[33]^r[26]^r[23]^r[22]^r[21]^r[20]^r[15]^r[14]^r[11]^r[7]^r[6]^r[5]^r[3]^r[2]^r[1]^g[240]^g[241]^g[246]^g[247]^g[248]^g[249]^g[250]^g[251]^g[254];
	g_next[243] = r[62]^r[58]^r[57]^r[54]^r[53]^r[52]^r[49]^r[48]^r[47]^r[44]^r[40]^r[39]^r[38]^r[36]^r[35]^r[32]^r[31]^r[29]^r[27]^r[26]^r[21]^r[20]^r[19]^r[17]^r[16]^r[14]^r[13]^r[8]^r[6]^r[0]^g[241]^g[242]^g[247]^g[248]^g[249]^g[250]^g[251]^g[252];
	g_next[244] = r[57]^r[52]^r[51]^r[49]^r[48]^r[47]^r[45]^r[38]^r[37]^r[33]^r[31]^r[29]^r[19]^r[18]^r[17]^r[15]^r[14]^r[13]^r[12]^r[11]^r[9]^r[8]^r[6]^r[3]^r[2]^g[242]^g[243]^g[248]^g[249]^g[250]^g[251]^g[252]^g[253];
	g_next[245] = r[62]^r[59]^r[53]^r[52]^r[50]^r[49]^r[48]^r[44]^r[39]^r[37]^r[36]^r[35]^r[34]^r[31]^r[28]^r[27]^r[23]^r[22]^r[18]^r[17]^r[16]^r[13]^r[11]^r[7]^r[6]^r[4]^r[3]^g[243]^g[244]^g[249]^g[250]^g[251]^g[252]^g[253]^g[254];
	g_next[246] = r[61]^r[59]^r[56]^r[51]^r[50]^r[49]^r[46]^r[45]^r[43]^r[42]^r[41]^r[39]^r[38]^r[37]^r[33]^r[30]^r[27]^r[26]^r[25]^r[23]^r[20]^r[18]^r[16]^r[15]^r[14]^r[12]^r[11]^r[10]^r[9]^r[8]^r[3]^r[2]^r[1]^g[240]^g[244]^g[245]^g[250]^g[251]^g[252]^g[253]^g[254];
	g_next[247] = r[57]^r[53]^r[51]^r[49]^r[46]^r[41]^r[38]^r[37]^r[35]^r[30]^r[28]^r[25]^r[22]^r[21]^r[20]^r[19]^r[18]^r[17]^r[16]^r[12]^r[11]^r[8]^r[7]^r[6]^r[4]^r[0]^g[241]^g[245]^g[246]^g[251]^g[252]^g[253]^g[254];
	g_next[248] = r[58]^r[57]^r[56]^r[53]^r[49]^r[46]^r[39]^r[37]^r[36]^r[33]^r[31]^r[28]^r[27]^r[25]^r[22]^r[21]^r[20]^r[19]^r[18]^r[17]^r[13]^r[10]^r[7]^r[6]^r[3]^r[2]^g[240]^g[242]^g[246]^g[247]^g[252]^g[253]^g[254];
	g_next[249] = r[60]^r[58]^r[56]^r[55]^r[51]^r[49]^r[47]^r[46]^r[45]^r[42]^r[41]^r[40]^r[38]^r[30]^r[29]^r[28]^r[26]^r[25]^r[24]^r[22]^r[19]^r[18]^r[16]^r[15]^r[12]^r[9]^r[5]^r[0]^g[241]^g[243]^g[247]^g[248]^g[253]^g[254];
	g_next[250] = r[61]^r[58]^r[56]^r[51]^r[50]^r[49]^r[47]^r[45]^r[43]^r[40]^r[38]^r[37]^r[35]^r[33]^r[30]^r[29]^r[26]^r[24]^r[22]^r[20]^r[19]^r[18]^r[12]^r[11]^r[7]^r[2]^g[240]^g[242]^g[244]^g[248]^g[249]^g[254];
	g_next[251] = r[60]^r[58]^r[57]^r[56]^r[52]^r[50]^r[49]^r[44]^r[42]^r[41]^r[40]^r[37]^r[35]^r[30]^r[29]^r[27]^r[25]^r[22]^r[21]^r[20]^r[18]^r[16]^r[15]^r[14]^r[13]^r[12]^r[11]^r[10]^r[8]^r[7]^r[6]^r[5]^r[0]^g[241]^g[243]^g[245]^g[249]^g[250];
	g_next[252] = r[59]^r[57]^r[56]^r[55]^r[54]^r[52]^r[46]^r[44]^r[41]^r[39]^r[36]^r[34]^r[28]^r[25]^r[23]^r[20]^r[19]^r[16]^r[14]^r[10]^r[8]^r[7]^r[6]^r[5]^r[4]^r[3]^g[242]^g[244]^g[246]^g[250]^g[251];
	g_next[253] = r[60]^r[56]^r[52]^r[50]^r[49]^r[46]^r[45]^r[44]^r[42]^r[39]^r[38]^r[37]^r[35]^r[34]^r[30]^r[29]^r[28]^r[27]^r[26]^r[25]^r[24]^r[23]^r[20]^r[16]^r[12]^r[11]^r[10]^r[9]^r[5]^r[2]^g[243]^g[245]^g[247]^g[251]^g[252];
	g_next[254] = r[56]^r[54]^r[51]^r[50]^r[49]^r[46]^r[45]^r[44]^r[43]^r[37]^r[36]^r[34]^r[27]^r[26]^r[25]^r[23]^r[20]^r[19]^r[18]^r[13]^r[12]^r[10]^r[9]^r[8]^r[7]^r[6]^r[5]^g[244]^g[246]^g[248]^g[252]^g[253];
	g_next[255] = r[63]^r[60]^r[57]^r[54]^r[51]^r[48]^r[46]^r[45]^r[44]^r[42]^r[40]^r[39]^r[38]^r[34]^r[33]^r[30]^r[29]^r[27]^r[25]^r[21]^r[17]^r[15]^r[13]^r[10]^r[6]^r[5]^r[3]^r[2]^r[0]^g[256]^g[258]^g[259]^g[262]^g[263]^g[267]^g[269];
	g_next[256] = r[60]^r[51]^r[50]^r[48]^r[44]^r[43]^r[39]^r[38]^r[37]^r[36]^r[31]^r[30]^r[27]^r[23]^r[22]^r[19]^r[15]^r[14]^r[12]^r[11]^r[10]^r[9]^r[0]^g[255]^g[256]^g[257]^g[258]^g[260]^g[262]^g[264]^g[267]^g[268]^g[269];
	g_next[257] = r[60]^r[57]^r[51]^r[50]^r[43]^r[42]^r[40]^r[36]^r[33]^r[32]^r[31]^r[28]^r[27]^r[26]^r[25]^r[24]^r[20]^r[19]^r[18]^r[13]^r[10]^g[256]^g[257]^g[258]^g[259]^g[261]^g[263]^g[265]^g[268]^g[269];
	g_next[258] = r[60]^r[58]^r[54]^r[52]^r[50]^r[46]^r[43]^r[42]^r[40]^r[39]^r[36]^r[32]^r[24]^r[23]^r[20]^r[16]^r[15]^r[14]^r[11]^r[9]^r[7]^r[6]^r[1]^g[255]^g[257]^g[258]^g[259]^g[260]^g[262]^g[264]^g[266]^g[269];
	g_next[259] = r[60]^r[57]^r[54]^r[52]^r[51]^r[50]^r[44]^r[43]^r[42]^r[38]^r[37]^r[28]^r[26]^r[24]^r[21]^r[20]^r[17]^r[15]^r[14]^r[12]^r[11]^r[7]^r[6]^r[4]^r[3]^g[256]^g[258]^g[259]^g[260]^g[261]^g[263]^g[265]^g[267];
	g_next[260] = r[62]^r[60]^r[59]^r[56]^r[53]^r[51]^r[47]^r[46]^r[43]^r[42]^r[41]^r[40]^r[39]^r[38]^r[37]^r[35]^r[32]^r[30]^r[29]^r[22]^r[17]^r[14]^r[11]^r[10]^r[9]^r[8]^r[7]^r[5]^r[4]^r[2]^g[257]^g[259]^g[260]^g[261]^g[262]^g[264]^g[266]^g[268];
	g_next[261] = r[60]^r[59]^r[57]^r[56]^r[52]^r[51]^r[50]^r[48]^r[47]^r[45]^r[44]^r[43]^r[40]^r[39]^r[38]^r[35]^r[32]^r[28]^r[26]^r[23]^r[21]^r[20]^r[18]^r[16]^r[15]^r[14]^r[11]^r[10]^r[8]^r[7]^r[5]^r[4]^r[1]^r[0]^g[258]^g[260]^g[261]^g[262]^g[263]^g[265]^g[267]^g[269];
	g_next[262] = r[62]^r[60]^r[58]^r[56]^r[54]^r[53]^r[52]^r[50]^r[48]^r[47]^r[46]^r[43]^r[42]^r[40]^r[34]^r[32]^r[31]^r[30]^r[29]^r[28]^r[26]^r[25]^r[22]^r[19]^r[15]^r[13]^r[12]^r[9]^r[8]^r[6]^r[5]^r[4]^r[0]^g[255]^g[259]^g[261]^g[262]^g[263]^g[264]^g[266]^g[268];
	g_next[263] = r[57]^r[53]^r[51]^r[50]^r[47]^r[45]^r[43]^r[41]^r[39]^r[37]^r[36]^r[31]^r[30]^r[29]^r[26]^r[23]^r[21]^r[19]^r[18]^r[15]^r[11]^r[9]^r[6]^r[5]^r[0]^g[255]^g[256]^g[260]^g[262]^g[263]^g[264]^g[265]^g[267]^g[269];
	g_next[264] = r[53]^r[51]^r[43]^r[39]^r[37]^r[36]^r[35]^r[32]^r[31]^r[30]^r[26]^r[24]^r[20]^r[18]^r[17]^r[16]^r[14]^r[13]^r[12]^r[11]^r[10]^r[9]^r[6]^r[5]^r[3]^r[2]^g[256]^g[257]^g[261]^g[263]^g[264]^g[265]^g[266]^g[268];
	g_next[265] = r[61]^r[58]^r[57]^r[55]^r[53]^r[52]^r[51]^r[50]^r[49]^r[46]^r[40]^r[37]^r[36]^r[35]^r[34]^r[29]^r[28]^r[23]^r[22]^r[21]^r[19]^r[16]^r[15]^r[14]^r[9]^r[7]^r[5]^r[4]^r[3]^r[1]^r[0]^g[257]^g[258]^g[262]^g[264]^g[265]^g[266]^g[267]^g[269];
	g_next[266] = r[58]^r[55]^r[53]^r[47]^r[46]^r[44]^r[41]^r[39]^r[38]^r[36]^r[34]^r[31]^r[23]^r[22]^r[17]^r[16]^r[15]^r[11]^r[9]^r[7]^r[5]^r[4]^r[2]^r[0]^g[255]^g[258]^g[259]^g[263]^g[265]^g[266]^g[267]^g[268];
	g_next[267] = r[58]^r[57]^r[53]^r[51]^r[50]^r[49]^r[47]^r[40]^r[38]^r[37]^r[36]^r[34]^r[33]^r[30]^r[27]^r[25]^r[24]^r[18]^r[16]^r[14]^r[13]^r[12]^r[11]^r[10]^r[9]^r[6]^r[5]^r[1]^g[255]^g[256]^g[259]^g[260]^g[264]^g[266]^g[267]^g[268]^g[269];
	g_next[268] = r[59]^r[58]^r[55]^r[52]^r[51]^r[47]^r[43]^r[40]^r[39]^r[37]^r[36]^r[35]^r[34]^r[31]^r[30]^r[29]^r[28]^r[27]^r[19]^r[18]^r[15]^r[13]^r[9]^r[8]^r[7]^r[6]^r[5]^r[3]^r[0]^g[256]^g[257]^g[260]^g[261]^g[265]^g[267]^g[268]^g[269];
	g_next[269] = r[61]^r[59]^r[57]^r[55]^r[53]^r[51]^r[50]^r[49]^r[47]^r[46]^r[45]^r[41]^r[39]^r[38]^r[36]^r[35]^r[34]^r[33]^r[28]^r[27]^r[24]^r[23]^r[21]^r[19]^r[18]^r[17]^r[16]^r[15]^r[14]^r[13]^r[10]^r[9]^r[7]^r[3]^r[2]^r[1]^g[255]^g[257]^g[258]^g[261]^g[262]^g[266]^g[268]^g[269];
	g_next[270] = r[63]^r[52]^r[48]^r[46]^r[42]^r[41]^r[36]^r[33]^r[32]^r[29]^r[24]^r[22]^r[21]^r[19]^r[14]^r[10]^r[9]^r[8]^r[3]^r[2]^r[1]^r[0]^g[271]^g[273]^g[274]^g[275]^g[276]^g[278]^g[279]^g[280]^g[282]^g[283];
	g_next[271] = r[57]^r[55]^r[52]^r[51]^r[50]^r[48]^r[45]^r[44]^r[42]^r[40]^r[38]^r[36]^r[35]^r[33]^r[32]^r[31]^r[26]^r[25]^r[24]^r[23]^r[20]^r[19]^r[17]^r[16]^r[14]^r[13]^r[10]^r[5]^r[4]^g[271]^g[272]^g[273]^g[277]^g[278]^g[281]^g[282]^g[284];
	g_next[272] = r[58]^r[57]^r[55]^r[52]^r[48]^r[47]^r[45]^r[44]^r[41]^r[39]^r[38]^r[37]^r[36]^r[35]^r[31]^r[30]^r[28]^r[27]^r[26]^r[23]^r[22]^r[21]^r[20]^r[19]^r[16]^r[14]^r[12]^r[9]^r[7]^r[5]^r[4]^r[3]^r[1]^g[270]^g[272]^g[273]^g[274]^g[278]^g[279]^g[282]^g[283];
	g_next[273] = r[61]^r[58]^r[57]^r[54]^r[53]^r[51]^r[50]^r[48]^r[42]^r[40]^r[36]^r[33]^r[30]^r[26]^r[25]^r[24]^r[23]^r[22]^r[20]^r[19]^r[18]^r[17]^r[16]^r[15]^r[9]^r[6]^r[0]^g[270]^g[271]^g[273]^g[274]^g[275]^g[279]^g[280]^g[283]^g[284];
	g_next[274] = r[61]^r[57]^r[56]^r[54]^r[52]^r[47]^r[44]^r[42]^r[41]^r[40]^r[38]^r[36]^r[32]^r[31]^r[28]^r[27]^r[26]^r[23]^r[22]^r[20]^r[17]^r[16]^r[14]^r[13]^r[12]^r[11]^r[10]^r[8]^r[7]^r[4]^r[2]^r[0]^g[271]^g[272]^g[274]^g[275]^g[276]^g[280]^g[281]^g[284];
	g_next[275] = r[58]^r[57]^r[52]^r[51]^r[50]^r[46]^r[45]^r[44]^r[43]^r[41]^r[39]^r[36]^r[34]^r[32]^r[25]^r[24]^r[23]^r[16]^r[14]^r[12]^r[11]^r[10]^r[8]^r[6]^r[5]^r[4]^r[2]^g[270]^g[272]^g[273]^g[275]^g[276]^g[277]^g[281]^g[282];
	g_next[276] = r[60]^r[59]^r[57]^r[54]^r[53]^r[48]^r[44]^r[42]^r[41]^r[40]^r[38]^r[37]^r[33]^r[30]^r[28]^r[26]^r[25]^r[23]^r[22]^r[21]^r[18]^r[17]^r[12]^r[11]^r[10]^r[9]^r[5]^r[3]^r[2]^r[0]^g[270]^g[271]^g[273]^g[274]^g[276]^g[277]^g[278]^g[282]^g[283];
	g_next[277] = r[62]^r[60]^r[57]^r[56]^r[52]^r[51]^r[48]^r[47]^r[46]^r[45]^r[44]^r[43]^r[42]^r[40]^r[32]^r[31]^r[28]^r[26]^r[25]^r[22]^r[20]^r[19]^r[15]^r[13]^r[12]^r[10]^r[9]^r[6]^r[5]^r[0]^g[270]^g[271]^g[272]^g[274]^g[275]^g[277]^g[278]^g[279]^g[283]^g[284];
	g_next[278] = r[60]^r[59]^r[57]^r[54]^r[49]^r[48]^r[47]^r[44]^r[43]^r[41]^r[40]^r[38]^r[34]^r[28]^r[26]^r[21]^r[20]^r[18]^r[17]^r[15]^r[12]^r[5]^r[4]^r[1]^r[0]^g[271]^g[272]^g[273]^g[275]^g[276]^g[278]^g[279]^g[280]^g[284];
	g_next[279] = r[62]^r[60]^r[58]^r[57]^r[48]^r[44]^r[43]^r[41]^r[40]^r[39]^r[36]^r[31]^r[30]^r[28]^r[27]^r[25]^r[24]^r[23]^r[21]^r[20]^r[19]^r[18]^r[17]^r[15]^r[14]^r[13]^r[12]^r[4]^r[3]^r[2]^r[1]^r[0]^g[270]^g[272]^g[273]^g[274]^g[276]^g[277]^g[279]^g[280]^g[281];
	g_next[280] = r[60]^r[57]^r[54]^r[53]^r[52]^r[51]^r[44]^r[43]^r[37]^r[34]^r[31]^r[30]^r[29]^r[21]^r[17]^r[14]^r[13]^r[12]^r[9]^r[8]^r[5]^r[4]^r[3]^g[270]^g[271]^g[273]^g[274]^g[275]^g[277]^g[278]^g[280]^g[281]^g[282];
	g_next[281] = r[60]^r[57]^r[55]^r[54]^r[53]^r[47]^r[44]^r[41]^r[39]^r[38]^r[36]^r[34]^r[31]^r[29]^r[20]^r[18]^r[16]^r[12]^r[10]^r[9]^r[8]^r[7]^r[4]^r[2]^r[1]^r[0]^g[270]^g[271]^g[272]^g[274]^g[275]^g[276]^g[278]^g[279]^g[281]^g[282]^g[283];
	g_next[282] = r[60]^r[53]^r[52]^r[51]^r[47]^r[45]^r[44]^r[43]^r[42]^r[41]^r[40]^r[39]^r[38]^r[33]^r[32]^r[31]^r[29]^r[25]^r[21]^r[19]^r[18]^r[17]^r[16]^r[14]^r[13]^r[11]^r[10]^r[9]^r[8]^r[7]^r[4]^r[3]^r[1]^g[270]^g[271]^g[272]^g[273]^g[275]^g[276]^g[277]^g[279]^g[280]^g[282]^g[283]^g[284];
	g_next[283] = r[60]^r[59]^r[58]^r[55]^r[52]^r[51]^r[47]^r[46]^r[36]^r[35]^r[32]^r[31]^r[30]^r[29]^r[26]^r[24]^r[20]^r[19]^r[17]^r[15]^r[13]^r[12]^r[8]^r[7]^r[6]^r[4]^r[3]^r[2]^g[271]^g[272]^g[273]^g[274]^g[276]^g[277]^g[278]^g[280]^g[281]^g[283]^g[284];
	g_next[284] = r[61]^r[59]^r[57]^r[55]^r[49]^r[47]^r[46]^r[41]^r[40]^r[39]^r[38]^r[35]^r[33]^r[30]^r[27]^r[25]^r[23]^r[22]^r[21]^r[19]^r[18]^r[15]^r[14]^r[13]^r[12]^r[10]^r[8]^r[7]^r[3]^r[1]^g[270]^g[272]^g[273]^g[274]^g[275]^g[277]^g[278]^g[279]^g[281]^g[282]^g[284];
	g_next[285] = r[63]^r[60]^r[58]^r[57]^r[54]^r[53]^r[52]^r[51]^r[50]^r[48]^r[45]^r[43]^r[41]^r[39]^r[38]^r[37]^r[36]^r[33]^r[32]^r[30]^r[27]^r[26]^r[23]^r[22]^r[20]^r[19]^r[15]^r[13]^r[12]^r[11]^r[9]^r[8]^r[6]^r[4]^r[3]^r[1]^r[0]^g[287]^g[289]^g[291]^g[292]^g[293]^g[295]^g[297]^g[299];
	g_next[286] = r[59]^r[58]^r[55]^r[54]^r[53]^r[52]^r[48]^r[45]^r[43]^r[42]^r[39]^r[38]^r[36]^r[35]^r[32]^r[31]^r[30]^r[27]^r[26]^r[25]^r[20]^r[19]^r[17]^r[16]^r[13]^r[12]^r[8]^r[5]^r[2]^r[0]^g[285]^g[287]^g[288]^g[289]^g[290]^g[291]^g[294]^g[295]^g[296]^g[297]^g[298]^g[299];
	g_next[287] = r[59]^r[52]^r[47]^r[46]^r[41]^r[39]^r[36]^r[35]^r[33]^r[32]^r[31]^r[28]^r[25]^r[23]^r[21]^r[19]^r[18]^r[17]^r[15]^r[12]^r[9]^r[7]^r[5]^r[4]^r[1]^g[286]^g[288]^g[289]^g[290]^g[291]^g[292]^g[295]^g[296]^g[297]^g[298]^g[299];
	g_next[288] = r[61]^r[56]^r[53]^r[51]^r[50]^r[45]^r[43]^r[42]^r[40]^r[39]^r[34]^r[31]^r[29]^r[28]^r[27]^r[26]^r[25]^r[24]^r[23]^r[22]^r[21]^r[20]^r[17]^r[15]^r[13]^r[12]^r[11]^r[7]^r[5]^r[4]^r[1]^r[0]^g[285]^g[287]^g[289]^g[290]^g[291]^g[292]^g[293]^g[296]^g[297]^g[298]^g[299];
	g_next[289] = r[61]^r[58]^r[56]^r[55]^r[53]^r[51]^r[48]^r[46]^r[45]^r[43]^r[42]^r[41]^r[40]^r[39]^r[38]^r[28]^r[27]^r[25]^r[23]^r[22]^r[21]^r[20]^r[19]^r[17]^r[13]^r[11]^r[9]^r[8]^r[5]^r[3]^r[2]^r[0]^g[286]^g[288]^g[290]^g[291]^g[292]^g[293]^g[294]^g[297]^g[298]^g[299];
	g_next[290] = r[60]^r[58]^r[52]^r[48]^r[45]^r[41]^r[40]^r[39]^r[38]^r[36]^r[33]^r[32]^r[31]^r[27]^r[26]^r[25]^r[23]^r[22]^r[21]^r[20]^r[19]^r[16]^r[15]^r[11]^r[8]^r[7]^r[6]^r[5]^r[4]^r[3]^r[2]^r[1]^r[0]^g[285]^g[287]^g[289]^g[291]^g[292]^g[293]^g[294]^g[295]^g[298]^g[299];
	g_next[291] = r[59]^r[56]^r[54]^r[52]^r[49]^r[48]^r[45]^r[44]^r[43]^r[41]^r[37]^r[34]^r[33]^r[31]^r[25]^r[24]^r[22]^r[19]^r[17]^r[16]^r[14]^r[12]^r[11]^r[10]^r[8]^r[7]^r[4]^r[3]^r[1]^r[0]^g[286]^g[288]^g[290]^g[292]^g[293]^g[294]^g[295]^g[296]^g[299];
	g_next[292] = r[61]^r[56]^r[51]^r[48]^r[45]^r[43]^r[42]^r[41]^r[40]^r[39]^r[34]^r[33]^r[31]^r[27]^r[25]^r[24]^r[22]^r[21]^r[20]^r[19]^r[18]^r[17]^r[15]^r[12]^r[11]^r[10]^r[8]^r[1]^g[285]^g[287]^g[289]^g[291]^g[293]^g[294]^g[295]^g[296]^g[297];
	g_next[293] = r[61]^r[59]^r[58]^r[54]^r[53]^r[51]^r[49]^r[47]^r[45]^r[44]^r[41]^r[40]^r[38]^r[34]^r[31]^r[29]^r[25]^r[24]^r[23]^r[20]^r[16]^r[14]^r[13]^r[11]^r[10]^r[1]^g[285]^g[286]^g[288]^g[290]^g[292]^g[294]^g[295]^g[296]^g[297]^g[298];
	g_next[294] = r[62]^r[58]^r[57]^r[54]^r[53]^r[51]^r[47]^r[46]^r[45]^r[44]^r[43]^r[42]^r[40]^r[39]^r[38]^r[37]^r[35]^r[34]^r[32]^r[31]^r[30]^r[28]^r[26]^r[22]^r[16]^r[15]^r[14]^r[12]^r[11]^r[10]^r[8]^r[7]^r[6]^r[5]^r[4]^r[3]^r[2]^g[285]^g[286]^g[287]^g[289]^g[291]^g[293]^g[295]^g[296]^g[297]^g[298]^g[299];
	g_next[295] = r[54]^r[52]^r[51]^r[48]^r[47]^r[45]^r[44]^r[43]^r[42]^r[41]^r[39]^r[37]^r[35]^r[34]^r[33]^r[32]^r[31]^r[30]^r[27]^r[24]^r[22]^r[20]^r[19]^r[17]^r[14]^r[13]^r[12]^r[11]^r[9]^r[7]^r[5]^r[2]^r[1]^g[286]^g[287]^g[288]^g[290]^g[292]^g[294]^g[296]^g[297]^g[298]^g[299];
	g_next[296] = r[62]^r[57]^r[54]^r[53]^r[52]^r[51]^r[48]^r[47]^r[45]^r[44]^r[42]^r[41]^r[40]^r[39]^r[37]^r[32]^r[31]^r[29]^r[25]^r[24]^r[22]^r[21]^r[20]^r[19]^r[16]^r[15]^r[14]^r[12]^r[11]^r[7]^r[5]^r[2]^r[1]^r[0]^g[285]^g[287]^g[288]^g[289]^g[291]^g[293]^g[295]^g[297]^g[298]^g[299];
	g_next[297] = r[60]^r[58]^r[57]^r[55]^r[54]^r[53]^r[51]^r[50]^r[49]^r[47]^r[39]^r[37]^r[35]^r[34]^r[33]^r[31]^r[29]^r[28]^r[27]^r[23]^r[22]^r[21]^r[20]^r[18]^r[15]^r[14]^r[10]^r[7]^r[6]^r[3]^r[1]^r[0]^g[286]^g[288]^g[289]^g[290]^g[292]^g[294]^g[296]^g[298]^g[299];
	g_next[298] = r[60]^r[58]^r[57]^r[55]^r[54]^r[52]^r[51]^r[50]^r[47]^r[46]^r[44]^r[42]^r[41]^r[39]^r[37]^r[35]^r[34]^r[32]^r[31]^r[30]^r[26]^r[21]^r[19]^r[17]^r[14]^r[12]^r[11]^r[10]^r[7]^r[6]^r[3]^r[2]^r[1]^r[0]^g[285]^g[287]^g[289]^g[290]^g[291]^g[293]^g[295]^g[297]^g[299];
	g_next[299] = r[60]^r[59]^r[57]^r[55]^r[52]^r[51]^r[50]^r[49]^r[47]^r[42]^r[41]^r[40]^r[37]^r[35]^r[33]^r[32]^r[31]^r[28]^r[27]^r[23]^r[18]^r[16]^r[15]^r[12]^r[11]^r[7]^r[5]^r[2]^r[1]^g[286]^g[288]^g[290]^g[291]^g[292]^g[294]^g[296]^g[298];
	return g_next;
endfunction

(* noinline *)
function Vector#(40, Bit#(15)) get_syndrome(Bit#(300) g);
	Vector#(40, Bit#(15)) syndrome = replicate(0);
	syndrome[0][0] = g[0];
	syndrome[0][1] = g[1];
	syndrome[0][2] = g[2];
	syndrome[0][3] = g[3];
	syndrome[0][4] = g[4];
	syndrome[0][5] = g[5];
	syndrome[0][6] = g[6];
	syndrome[0][7] = g[7];
	syndrome[0][8] = g[8];
	syndrome[0][9] = g[9];
	syndrome[0][10] = g[10];
	syndrome[0][11] = g[11];
	syndrome[0][12] = g[12];
	syndrome[0][13] = g[13];
	syndrome[0][14] = g[14];
	syndrome[1][0] = g[0];
	syndrome[1][1] = g[8];
	syndrome[1][2] = g[1]^g[8];
	syndrome[1][3] = g[9];
	syndrome[1][4] = g[2]^g[9];
	syndrome[1][5] = g[10];
	syndrome[1][6] = g[3]^g[10];
	syndrome[1][7] = g[11];
	syndrome[1][8] = g[4]^g[11];
	syndrome[1][9] = g[12];
	syndrome[1][10] = g[5]^g[12];
	syndrome[1][11] = g[13];
	syndrome[1][12] = g[6]^g[13];
	syndrome[1][13] = g[14];
	syndrome[1][14] = g[7]^g[14];
	syndrome[2][0] = g[15];
	syndrome[2][1] = g[16];
	syndrome[2][2] = g[17];
	syndrome[2][3] = g[18];
	syndrome[2][4] = g[19];
	syndrome[2][5] = g[20];
	syndrome[2][6] = g[21];
	syndrome[2][7] = g[22];
	syndrome[2][8] = g[23];
	syndrome[2][9] = g[24];
	syndrome[2][10] = g[25];
	syndrome[2][11] = g[26];
	syndrome[2][12] = g[27];
	syndrome[2][13] = g[28];
	syndrome[2][14] = g[29];
	syndrome[3][0] = g[0];
	syndrome[3][1] = g[4]^g[11];
	syndrome[3][2] = g[4]^g[8]^g[11];
	syndrome[3][3] = g[12];
	syndrome[3][4] = g[1]^g[8]^g[12];
	syndrome[3][5] = g[5]^g[12];
	syndrome[3][6] = g[5]^g[9]^g[12];
	syndrome[3][7] = g[13];
	syndrome[3][8] = g[2]^g[9]^g[13];
	syndrome[3][9] = g[6]^g[13];
	syndrome[3][10] = g[6]^g[10]^g[13];
	syndrome[3][11] = g[14];
	syndrome[3][12] = g[3]^g[10]^g[14];
	syndrome[3][13] = g[7]^g[14];
	syndrome[3][14] = g[7]^g[11]^g[14];
	syndrome[4][0] = g[30];
	syndrome[4][1] = g[31];
	syndrome[4][2] = g[32];
	syndrome[4][3] = g[33];
	syndrome[4][4] = g[34];
	syndrome[4][5] = g[35];
	syndrome[4][6] = g[36];
	syndrome[4][7] = g[37];
	syndrome[4][8] = g[38];
	syndrome[4][9] = g[39];
	syndrome[4][10] = g[40];
	syndrome[4][11] = g[41];
	syndrome[4][12] = g[42];
	syndrome[4][13] = g[43];
	syndrome[4][14] = g[44];
	syndrome[5][0] = g[15];
	syndrome[5][1] = g[23];
	syndrome[5][2] = g[16]^g[23];
	syndrome[5][3] = g[24];
	syndrome[5][4] = g[17]^g[24];
	syndrome[5][5] = g[25];
	syndrome[5][6] = g[18]^g[25];
	syndrome[5][7] = g[26];
	syndrome[5][8] = g[19]^g[26];
	syndrome[5][9] = g[27];
	syndrome[5][10] = g[20]^g[27];
	syndrome[5][11] = g[28];
	syndrome[5][12] = g[21]^g[28];
	syndrome[5][13] = g[29];
	syndrome[5][14] = g[22]^g[29];
	syndrome[6][0] = g[45];
	syndrome[6][1] = g[46];
	syndrome[6][2] = g[47];
	syndrome[6][3] = g[48];
	syndrome[6][4] = g[49];
	syndrome[6][5] = g[50];
	syndrome[6][6] = g[51];
	syndrome[6][7] = g[52];
	syndrome[6][8] = g[53];
	syndrome[6][9] = g[54];
	syndrome[6][10] = g[55];
	syndrome[6][11] = g[56];
	syndrome[6][12] = g[57];
	syndrome[6][13] = g[58];
	syndrome[6][14] = g[59];
	syndrome[7][0] = g[0];
	syndrome[7][1] = g[2]^g[9]^g[13];
	syndrome[7][2] = g[2]^g[4]^g[9]^g[11]^g[13];
	syndrome[7][3] = g[6]^g[13];
	syndrome[7][4] = g[4]^g[6]^g[8]^g[11]^g[13];
	syndrome[7][5] = g[6]^g[10]^g[13];
	syndrome[7][6] = g[6]^g[10]^g[12]^g[13];
	syndrome[7][7] = g[14];
	syndrome[7][8] = g[1]^g[8]^g[12]^g[14];
	syndrome[7][9] = g[3]^g[10]^g[14];
	syndrome[7][10] = g[3]^g[5]^g[10]^g[12]^g[14];
	syndrome[7][11] = g[7]^g[14];
	syndrome[7][12] = g[5]^g[7]^g[9]^g[12]^g[14];
	syndrome[7][13] = g[7]^g[11]^g[14];
	syndrome[7][14] = g[7]^g[11]^g[13]^g[14];
	syndrome[8][0] = g[60];
	syndrome[8][1] = g[61];
	syndrome[8][2] = g[62];
	syndrome[8][3] = g[63];
	syndrome[8][4] = g[64];
	syndrome[8][5] = g[65];
	syndrome[8][6] = g[66];
	syndrome[8][7] = g[67];
	syndrome[8][8] = g[68];
	syndrome[8][9] = g[69];
	syndrome[8][10] = g[70];
	syndrome[8][11] = g[71];
	syndrome[8][12] = g[72];
	syndrome[8][13] = g[73];
	syndrome[8][14] = g[74];
	syndrome[9][0] = g[30];
	syndrome[9][1] = g[38];
	syndrome[9][2] = g[31]^g[38];
	syndrome[9][3] = g[39];
	syndrome[9][4] = g[32]^g[39];
	syndrome[9][5] = g[40];
	syndrome[9][6] = g[33]^g[40];
	syndrome[9][7] = g[41];
	syndrome[9][8] = g[34]^g[41];
	syndrome[9][9] = g[42];
	syndrome[9][10] = g[35]^g[42];
	syndrome[9][11] = g[43];
	syndrome[9][12] = g[36]^g[43];
	syndrome[9][13] = g[44];
	syndrome[9][14] = g[37]^g[44];
	syndrome[10][0] = g[75];
	syndrome[10][1] = g[76];
	syndrome[10][2] = g[77];
	syndrome[10][3] = g[78];
	syndrome[10][4] = g[79];
	syndrome[10][5] = g[80];
	syndrome[10][6] = g[81];
	syndrome[10][7] = g[82];
	syndrome[10][8] = g[83];
	syndrome[10][9] = g[84];
	syndrome[10][10] = g[85];
	syndrome[10][11] = g[86];
	syndrome[10][12] = g[87];
	syndrome[10][13] = g[88];
	syndrome[10][14] = g[89];
	syndrome[11][0] = g[15];
	syndrome[11][1] = g[19]^g[26];
	syndrome[11][2] = g[19]^g[23]^g[26];
	syndrome[11][3] = g[27];
	syndrome[11][4] = g[16]^g[23]^g[27];
	syndrome[11][5] = g[20]^g[27];
	syndrome[11][6] = g[20]^g[24]^g[27];
	syndrome[11][7] = g[28];
	syndrome[11][8] = g[17]^g[24]^g[28];
	syndrome[11][9] = g[21]^g[28];
	syndrome[11][10] = g[21]^g[25]^g[28];
	syndrome[11][11] = g[29];
	syndrome[11][12] = g[18]^g[25]^g[29];
	syndrome[11][13] = g[22]^g[29];
	syndrome[11][14] = g[22]^g[26]^g[29];
	syndrome[12][0] = g[90];
	syndrome[12][1] = g[91];
	syndrome[12][2] = g[92];
	syndrome[12][3] = g[93];
	syndrome[12][4] = g[94];
	syndrome[12][5] = g[95];
	syndrome[12][6] = g[96];
	syndrome[12][7] = g[97];
	syndrome[12][8] = g[98];
	syndrome[12][9] = g[99];
	syndrome[12][10] = g[100];
	syndrome[12][11] = g[101];
	syndrome[12][12] = g[102];
	syndrome[12][13] = g[103];
	syndrome[12][14] = g[104];
	syndrome[13][0] = g[45];
	syndrome[13][1] = g[53];
	syndrome[13][2] = g[46]^g[53];
	syndrome[13][3] = g[54];
	syndrome[13][4] = g[47]^g[54];
	syndrome[13][5] = g[55];
	syndrome[13][6] = g[48]^g[55];
	syndrome[13][7] = g[56];
	syndrome[13][8] = g[49]^g[56];
	syndrome[13][9] = g[57];
	syndrome[13][10] = g[50]^g[57];
	syndrome[13][11] = g[58];
	syndrome[13][12] = g[51]^g[58];
	syndrome[13][13] = g[59];
	syndrome[13][14] = g[52]^g[59];
	syndrome[14][0] = g[105];
	syndrome[14][1] = g[106];
	syndrome[14][2] = g[107];
	syndrome[14][3] = g[108];
	syndrome[14][4] = g[109];
	syndrome[14][5] = g[110];
	syndrome[14][6] = g[111];
	syndrome[14][7] = g[112];
	syndrome[14][8] = g[113];
	syndrome[14][9] = g[114];
	syndrome[14][10] = g[115];
	syndrome[14][11] = g[116];
	syndrome[14][12] = g[117];
	syndrome[14][13] = g[118];
	syndrome[14][14] = g[119];
	syndrome[15][0] = g[0];
	syndrome[15][1] = g[1]^g[8]^g[12]^g[14];
	syndrome[15][2] = g[1]^g[2]^g[8]^g[9]^g[12]^g[13]^g[14];
	syndrome[15][3] = g[3]^g[10]^g[14];
	syndrome[15][4] = g[2]^g[3]^g[4]^g[9]^g[10]^g[11]^g[13]^g[14];
	syndrome[15][5] = g[3]^g[5]^g[10]^g[12]^g[14];
	syndrome[15][6] = g[3]^g[5]^g[6]^g[10]^g[12]^g[13]^g[14];
	syndrome[15][7] = g[7]^g[14];
	syndrome[15][8] = g[4]^g[6]^g[7]^g[8]^g[11]^g[13]^g[14];
	syndrome[15][9] = g[5]^g[7]^g[9]^g[12]^g[14];
	syndrome[15][10] = g[5]^g[6]^g[7]^g[9]^g[10]^g[12]^g[13]^g[14];
	syndrome[15][11] = g[7]^g[11]^g[14];
	syndrome[15][12] = g[6]^g[7]^g[10]^g[11]^g[12]^g[13]^g[14];
	syndrome[15][13] = g[7]^g[11]^g[13]^g[14];
	syndrome[15][14] = g[7]^g[11]^g[13];
	syndrome[16][0] = g[120];
	syndrome[16][1] = g[121];
	syndrome[16][2] = g[122];
	syndrome[16][3] = g[123];
	syndrome[16][4] = g[124];
	syndrome[16][5] = g[125];
	syndrome[16][6] = g[126];
	syndrome[16][7] = g[127];
	syndrome[16][8] = g[128];
	syndrome[16][9] = g[129];
	syndrome[16][10] = g[130];
	syndrome[16][11] = g[131];
	syndrome[16][12] = g[132];
	syndrome[16][13] = g[133];
	syndrome[16][14] = g[134];
	syndrome[17][0] = g[60];
	syndrome[17][1] = g[68];
	syndrome[17][2] = g[61]^g[68];
	syndrome[17][3] = g[69];
	syndrome[17][4] = g[62]^g[69];
	syndrome[17][5] = g[70];
	syndrome[17][6] = g[63]^g[70];
	syndrome[17][7] = g[71];
	syndrome[17][8] = g[64]^g[71];
	syndrome[17][9] = g[72];
	syndrome[17][10] = g[65]^g[72];
	syndrome[17][11] = g[73];
	syndrome[17][12] = g[66]^g[73];
	syndrome[17][13] = g[74];
	syndrome[17][14] = g[67]^g[74];
	syndrome[18][0] = g[135];
	syndrome[18][1] = g[136];
	syndrome[18][2] = g[137];
	syndrome[18][3] = g[138];
	syndrome[18][4] = g[139];
	syndrome[18][5] = g[140];
	syndrome[18][6] = g[141];
	syndrome[18][7] = g[142];
	syndrome[18][8] = g[143];
	syndrome[18][9] = g[144];
	syndrome[18][10] = g[145];
	syndrome[18][11] = g[146];
	syndrome[18][12] = g[147];
	syndrome[18][13] = g[148];
	syndrome[18][14] = g[149];
	syndrome[19][0] = g[30];
	syndrome[19][1] = g[34]^g[41];
	syndrome[19][2] = g[34]^g[38]^g[41];
	syndrome[19][3] = g[42];
	syndrome[19][4] = g[31]^g[38]^g[42];
	syndrome[19][5] = g[35]^g[42];
	syndrome[19][6] = g[35]^g[39]^g[42];
	syndrome[19][7] = g[43];
	syndrome[19][8] = g[32]^g[39]^g[43];
	syndrome[19][9] = g[36]^g[43];
	syndrome[19][10] = g[36]^g[40]^g[43];
	syndrome[19][11] = g[44];
	syndrome[19][12] = g[33]^g[40]^g[44];
	syndrome[19][13] = g[37]^g[44];
	syndrome[19][14] = g[37]^g[41]^g[44];
	syndrome[20][0] = g[150];
	syndrome[20][1] = g[151];
	syndrome[20][2] = g[152];
	syndrome[20][3] = g[153];
	syndrome[20][4] = g[154];
	syndrome[20][5] = g[155];
	syndrome[20][6] = g[156];
	syndrome[20][7] = g[157];
	syndrome[20][8] = g[158];
	syndrome[20][9] = g[159];
	syndrome[20][10] = g[160];
	syndrome[20][11] = g[161];
	syndrome[20][12] = g[162];
	syndrome[20][13] = g[163];
	syndrome[20][14] = g[164];
	syndrome[21][0] = g[75];
	syndrome[21][1] = g[83];
	syndrome[21][2] = g[76]^g[83];
	syndrome[21][3] = g[84];
	syndrome[21][4] = g[77]^g[84];
	syndrome[21][5] = g[85];
	syndrome[21][6] = g[78]^g[85];
	syndrome[21][7] = g[86];
	syndrome[21][8] = g[79]^g[86];
	syndrome[21][9] = g[87];
	syndrome[21][10] = g[80]^g[87];
	syndrome[21][11] = g[88];
	syndrome[21][12] = g[81]^g[88];
	syndrome[21][13] = g[89];
	syndrome[21][14] = g[82]^g[89];
	syndrome[22][0] = g[165];
	syndrome[22][1] = g[166];
	syndrome[22][2] = g[167];
	syndrome[22][3] = g[168];
	syndrome[22][4] = g[169];
	syndrome[22][5] = g[170];
	syndrome[22][6] = g[171];
	syndrome[22][7] = g[172];
	syndrome[22][8] = g[173];
	syndrome[22][9] = g[174];
	syndrome[22][10] = g[175];
	syndrome[22][11] = g[176];
	syndrome[22][12] = g[177];
	syndrome[22][13] = g[178];
	syndrome[22][14] = g[179];
	syndrome[23][0] = g[15];
	syndrome[23][1] = g[17]^g[24]^g[28];
	syndrome[23][2] = g[17]^g[19]^g[24]^g[26]^g[28];
	syndrome[23][3] = g[21]^g[28];
	syndrome[23][4] = g[19]^g[21]^g[23]^g[26]^g[28];
	syndrome[23][5] = g[21]^g[25]^g[28];
	syndrome[23][6] = g[21]^g[25]^g[27]^g[28];
	syndrome[23][7] = g[29];
	syndrome[23][8] = g[16]^g[23]^g[27]^g[29];
	syndrome[23][9] = g[18]^g[25]^g[29];
	syndrome[23][10] = g[18]^g[20]^g[25]^g[27]^g[29];
	syndrome[23][11] = g[22]^g[29];
	syndrome[23][12] = g[20]^g[22]^g[24]^g[27]^g[29];
	syndrome[23][13] = g[22]^g[26]^g[29];
	syndrome[23][14] = g[22]^g[26]^g[28]^g[29];
	syndrome[24][0] = g[180];
	syndrome[24][1] = g[181];
	syndrome[24][2] = g[182];
	syndrome[24][3] = g[183];
	syndrome[24][4] = g[184];
	syndrome[24][5] = g[185];
	syndrome[24][6] = g[186];
	syndrome[24][7] = g[187];
	syndrome[24][8] = g[188];
	syndrome[24][9] = g[189];
	syndrome[24][10] = g[190];
	syndrome[24][11] = g[191];
	syndrome[24][12] = g[192];
	syndrome[24][13] = g[193];
	syndrome[24][14] = g[194];
	syndrome[25][0] = g[90];
	syndrome[25][1] = g[98];
	syndrome[25][2] = g[91]^g[98];
	syndrome[25][3] = g[99];
	syndrome[25][4] = g[92]^g[99];
	syndrome[25][5] = g[100];
	syndrome[25][6] = g[93]^g[100];
	syndrome[25][7] = g[101];
	syndrome[25][8] = g[94]^g[101];
	syndrome[25][9] = g[102];
	syndrome[25][10] = g[95]^g[102];
	syndrome[25][11] = g[103];
	syndrome[25][12] = g[96]^g[103];
	syndrome[25][13] = g[104];
	syndrome[25][14] = g[97]^g[104];
	syndrome[26][0] = g[195];
	syndrome[26][1] = g[196];
	syndrome[26][2] = g[197];
	syndrome[26][3] = g[198];
	syndrome[26][4] = g[199];
	syndrome[26][5] = g[200];
	syndrome[26][6] = g[201];
	syndrome[26][7] = g[202];
	syndrome[26][8] = g[203];
	syndrome[26][9] = g[204];
	syndrome[26][10] = g[205];
	syndrome[26][11] = g[206];
	syndrome[26][12] = g[207];
	syndrome[26][13] = g[208];
	syndrome[26][14] = g[209];
	syndrome[27][0] = g[45];
	syndrome[27][1] = g[49]^g[56];
	syndrome[27][2] = g[49]^g[53]^g[56];
	syndrome[27][3] = g[57];
	syndrome[27][4] = g[46]^g[53]^g[57];
	syndrome[27][5] = g[50]^g[57];
	syndrome[27][6] = g[50]^g[54]^g[57];
	syndrome[27][7] = g[58];
	syndrome[27][8] = g[47]^g[54]^g[58];
	syndrome[27][9] = g[51]^g[58];
	syndrome[27][10] = g[51]^g[55]^g[58];
	syndrome[27][11] = g[59];
	syndrome[27][12] = g[48]^g[55]^g[59];
	syndrome[27][13] = g[52]^g[59];
	syndrome[27][14] = g[52]^g[56]^g[59];
	syndrome[28][0] = g[210];
	syndrome[28][1] = g[211];
	syndrome[28][2] = g[212];
	syndrome[28][3] = g[213];
	syndrome[28][4] = g[214];
	syndrome[28][5] = g[215];
	syndrome[28][6] = g[216];
	syndrome[28][7] = g[217];
	syndrome[28][8] = g[218];
	syndrome[28][9] = g[219];
	syndrome[28][10] = g[220];
	syndrome[28][11] = g[221];
	syndrome[28][12] = g[222];
	syndrome[28][13] = g[223];
	syndrome[28][14] = g[224];
	syndrome[29][0] = g[105];
	syndrome[29][1] = g[113];
	syndrome[29][2] = g[106]^g[113];
	syndrome[29][3] = g[114];
	syndrome[29][4] = g[107]^g[114];
	syndrome[29][5] = g[115];
	syndrome[29][6] = g[108]^g[115];
	syndrome[29][7] = g[116];
	syndrome[29][8] = g[109]^g[116];
	syndrome[29][9] = g[117];
	syndrome[29][10] = g[110]^g[117];
	syndrome[29][11] = g[118];
	syndrome[29][12] = g[111]^g[118];
	syndrome[29][13] = g[119];
	syndrome[29][14] = g[112]^g[119];
	syndrome[30][0] = g[225];
	syndrome[30][1] = g[226];
	syndrome[30][2] = g[227];
	syndrome[30][3] = g[228];
	syndrome[30][4] = g[229];
	syndrome[30][5] = g[230];
	syndrome[30][6] = g[231];
	syndrome[30][7] = g[232];
	syndrome[30][8] = g[233];
	syndrome[30][9] = g[234];
	syndrome[30][10] = g[235];
	syndrome[30][11] = g[236];
	syndrome[30][12] = g[237];
	syndrome[30][13] = g[238];
	syndrome[30][14] = g[239];
	syndrome[31][0] = g[0];
	syndrome[31][1] = g[4]^g[6]^g[7]^g[8]^g[11]^g[13]^g[14];
	syndrome[31][2] = g[1]^g[4]^g[6]^g[7]^g[11]^g[12]^g[13];
	syndrome[31][3] = g[5]^g[7]^g[9]^g[12]^g[14];
	syndrome[31][4] = g[1]^g[2]^g[5]^g[7]^g[8]^g[13];
	syndrome[31][5] = g[5]^g[6]^g[7]^g[9]^g[10]^g[12]^g[13]^g[14];
	syndrome[31][6] = g[3]^g[5]^g[6]^g[7]^g[9]^g[12]^g[13];
	syndrome[31][7] = g[7]^g[11]^g[14];
	syndrome[31][8] = g[2]^g[3]^g[4]^g[7]^g[9]^g[10]^g[13];
	syndrome[31][9] = g[6]^g[7]^g[10]^g[11]^g[12]^g[13]^g[14];
	syndrome[31][10] = g[3]^g[5]^g[6]^g[7]^g[11]^g[13];
	syndrome[31][11] = g[7]^g[11]^g[13]^g[14];
	syndrome[31][12] = g[3]^g[5]^g[6]^g[7]^g[10]^g[11]^g[12];
	syndrome[31][13] = g[7]^g[11]^g[13];
	syndrome[31][14] = g[11]^g[13]^g[14];
	syndrome[32][0] = g[240];
	syndrome[32][1] = g[241];
	syndrome[32][2] = g[242];
	syndrome[32][3] = g[243];
	syndrome[32][4] = g[244];
	syndrome[32][5] = g[245];
	syndrome[32][6] = g[246];
	syndrome[32][7] = g[247];
	syndrome[32][8] = g[248];
	syndrome[32][9] = g[249];
	syndrome[32][10] = g[250];
	syndrome[32][11] = g[251];
	syndrome[32][12] = g[252];
	syndrome[32][13] = g[253];
	syndrome[32][14] = g[254];
	syndrome[33][0] = g[120];
	syndrome[33][1] = g[128];
	syndrome[33][2] = g[121]^g[128];
	syndrome[33][3] = g[129];
	syndrome[33][4] = g[122]^g[129];
	syndrome[33][5] = g[130];
	syndrome[33][6] = g[123]^g[130];
	syndrome[33][7] = g[131];
	syndrome[33][8] = g[124]^g[131];
	syndrome[33][9] = g[132];
	syndrome[33][10] = g[125]^g[132];
	syndrome[33][11] = g[133];
	syndrome[33][12] = g[126]^g[133];
	syndrome[33][13] = g[134];
	syndrome[33][14] = g[127]^g[134];
	syndrome[34][0] = g[255];
	syndrome[34][1] = g[256];
	syndrome[34][2] = g[257];
	syndrome[34][3] = g[258];
	syndrome[34][4] = g[259];
	syndrome[34][5] = g[260];
	syndrome[34][6] = g[261];
	syndrome[34][7] = g[262];
	syndrome[34][8] = g[263];
	syndrome[34][9] = g[264];
	syndrome[34][10] = g[265];
	syndrome[34][11] = g[266];
	syndrome[34][12] = g[267];
	syndrome[34][13] = g[268];
	syndrome[34][14] = g[269];
	syndrome[35][0] = g[60];
	syndrome[35][1] = g[64]^g[71];
	syndrome[35][2] = g[64]^g[68]^g[71];
	syndrome[35][3] = g[72];
	syndrome[35][4] = g[61]^g[68]^g[72];
	syndrome[35][5] = g[65]^g[72];
	syndrome[35][6] = g[65]^g[69]^g[72];
	syndrome[35][7] = g[73];
	syndrome[35][8] = g[62]^g[69]^g[73];
	syndrome[35][9] = g[66]^g[73];
	syndrome[35][10] = g[66]^g[70]^g[73];
	syndrome[35][11] = g[74];
	syndrome[35][12] = g[63]^g[70]^g[74];
	syndrome[35][13] = g[67]^g[74];
	syndrome[35][14] = g[67]^g[71]^g[74];
	syndrome[36][0] = g[270];
	syndrome[36][1] = g[271];
	syndrome[36][2] = g[272];
	syndrome[36][3] = g[273];
	syndrome[36][4] = g[274];
	syndrome[36][5] = g[275];
	syndrome[36][6] = g[276];
	syndrome[36][7] = g[277];
	syndrome[36][8] = g[278];
	syndrome[36][9] = g[279];
	syndrome[36][10] = g[280];
	syndrome[36][11] = g[281];
	syndrome[36][12] = g[282];
	syndrome[36][13] = g[283];
	syndrome[36][14] = g[284];
	syndrome[37][0] = g[135];
	syndrome[37][1] = g[143];
	syndrome[37][2] = g[136]^g[143];
	syndrome[37][3] = g[144];
	syndrome[37][4] = g[137]^g[144];
	syndrome[37][5] = g[145];
	syndrome[37][6] = g[138]^g[145];
	syndrome[37][7] = g[146];
	syndrome[37][8] = g[139]^g[146];
	syndrome[37][9] = g[147];
	syndrome[37][10] = g[140]^g[147];
	syndrome[37][11] = g[148];
	syndrome[37][12] = g[141]^g[148];
	syndrome[37][13] = g[149];
	syndrome[37][14] = g[142]^g[149];
	syndrome[38][0] = g[285];
	syndrome[38][1] = g[286];
	syndrome[38][2] = g[287];
	syndrome[38][3] = g[288];
	syndrome[38][4] = g[289];
	syndrome[38][5] = g[290];
	syndrome[38][6] = g[291];
	syndrome[38][7] = g[292];
	syndrome[38][8] = g[293];
	syndrome[38][9] = g[294];
	syndrome[38][10] = g[295];
	syndrome[38][11] = g[296];
	syndrome[38][12] = g[297];
	syndrome[38][13] = g[298];
	syndrome[38][14] = g[299];
	syndrome[39][0] = g[30];
	syndrome[39][1] = g[32]^g[39]^g[43];
	syndrome[39][2] = g[32]^g[34]^g[39]^g[41]^g[43];
	syndrome[39][3] = g[36]^g[43];
	syndrome[39][4] = g[34]^g[36]^g[38]^g[41]^g[43];
	syndrome[39][5] = g[36]^g[40]^g[43];
	syndrome[39][6] = g[36]^g[40]^g[42]^g[43];
	syndrome[39][7] = g[44];
	syndrome[39][8] = g[31]^g[38]^g[42]^g[44];
	syndrome[39][9] = g[33]^g[40]^g[44];
	syndrome[39][10] = g[33]^g[35]^g[40]^g[42]^g[44];
	syndrome[39][11] = g[37]^g[44];
	syndrome[39][12] = g[35]^g[37]^g[39]^g[42]^g[44];
	syndrome[39][13] = g[37]^g[41]^g[44];
	syndrome[39][14] = g[37]^g[41]^g[43]^g[44];
	return syndrome;
endfunction
