function SubcodeInstruction page_0_get_instruction(UInt#(6) instr_counter);
	SubcodeInstruction ci;
	ci.offset = 0;
	ci.instructionVector = replicate(R1N256);
	case (instr_counter)
		6'd0 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd1 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd2 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd3 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd4 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd5 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd6 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd7 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = ML2N16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = R1N8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPR04N8; ci.instructionVector[10] = R0N8; end
		6'd8 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd9 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd10 : begin ci.offset = 60; ci.instructionVector[0] = ML2N16; end
		6'd11 : begin ci.offset = 30; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = ML2N8; ci.instructionVector[9] = SPCN8; ci.instructionVector[10] = SPCN16; end
		6'd12 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd13 : begin ci.offset = 24; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R1N16; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = ML2N16; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = R0N16; end
		6'd14 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = ML2N8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = ML2N16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = ML2R04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = R0N16; end
		6'd15 : begin ci.offset = 4; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = R0N8; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = ML2R04N8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = R0N32; ci.instructionVector[15] = R0N64; end
		6'd16 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd17 : begin ci.offset = 62; ci.instructionVector[0] = R14SPCN8; end
		6'd18 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd19 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = ML2N8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = ML2N16; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = R0N16; end
		6'd20 : begin ci.offset = 52; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = ML2R04N8; end
		6'd21 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = ML2N16; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = R1N8; ci.instructionVector[8] = R14SPCN8; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = R0N8; ci.instructionVector[13] = REPN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = ML2R04N8; ci.instructionVector[16] = R0N8; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; end
		6'd22 : begin ci.offset = 12; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = R1N8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = ML2R04N8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = R14SPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N32; end
		6'd23 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = ML2N8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = ML2R04N8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd24 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = ML2N16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; end
		6'd25 : begin ci.offset = 14; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPR04N8; ci.instructionVector[11] = ML2N8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N32; end
		6'd26 : begin ci.offset = 8; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = ML2R04N8; ci.instructionVector[6] = R14SPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = ML2N16; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = R0N16; ci.instructionVector[15] = REPR04N8; ci.instructionVector[16] = R0N8; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = R0N32; end
		6'd27 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = ML2R04N8; ci.instructionVector[5] = R0N8; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd28 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = ML2N16; ci.instructionVector[2] = R14SPCN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = R1N8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPR04N8; ci.instructionVector[9] = R0N8; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd29 : begin ci.offset = 0; ci.instructionVector[0] = ML2N8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = R0N64; ci.instructionVector[6] = R0N128; end
		6'd30 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd31 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd32 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd33 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd34 : begin ci.offset = 52; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPR04N8; end
		6'd35 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = ML2N8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = ML2N16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPR04N8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N16; end
		6'd36 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; end
		6'd37 : begin ci.offset = 12; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = R1N8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = ML2R04N8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = R14SPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N32; end
		6'd38 : begin ci.offset = 12; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = ML2N8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = R0N16; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = R0N32; end
		6'd39 : begin ci.offset = 2; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = R0N8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = R0N32; ci.instructionVector[12] = R0N64; end
		6'd40 : begin ci.offset = 28; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = REPR04N8; ci.instructionVector[10] = SPCN16; end
		6'd41 : begin ci.offset = 8; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = R14SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = ML2R04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd42 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = ML2N16; ci.instructionVector[2] = R14SPCN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = R1N8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPR04N8; ci.instructionVector[9] = R0N8; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = ML2R04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd43 : begin ci.offset = 0; ci.instructionVector[0] = ML2N8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = R0N64; ci.instructionVector[6] = R0N128; end
		6'd44 : begin ci.offset = 6; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = SPCN16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd45 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = R0N8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd46 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd47 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd48 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = ML2N8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = R14SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = R0N16; end
		6'd49 : begin ci.offset = 4; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = ML2R04N8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = R0N64; end
		6'd50 : begin ci.offset = 4; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = ML2N8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd51 : begin ci.offset = 0; ci.instructionVector[0] = REPR04N8; ci.instructionVector[1] = R0N8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd52 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = ML2N8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = ML2R04N8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd53 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd54 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd55 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd56 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = ML2R04N8; ci.instructionVector[5] = R0N8; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd57 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd58 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd59 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd60 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd61 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd62 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd63 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
	endcase
	return ci;
endfunction

function Codeword page_0_get_msg_bit_ind(UInt#(6) subcodeword_counter);
	Codeword msg_bit_ind=case (subcodeword_counter)
		6'd0: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd3: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd4: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd5: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd6: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd7: 256'b0000000000000111000101110111111100010111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd8: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd9: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd10: 256'b0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd11: 256'b0000000000000001000000010011111100000111011111110111111111111111000101110111111111111111111111111111111111111111111111111111111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd12: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd13: 256'b0000000000000000000000010001011100000001000101110011111111111111000000010111111101111111111111110111111111111111111111111111111100010111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd14: 256'b0000000000000000000000000000001100000000000101110001011101111111000000010001011100011111111111110011111111111111111111111111111100000001001111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd15: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001011100000000000000000000000000000001000000000000000100000011011111110000000000000111000101110111111100010111011111111111111111111111;
		6'd16: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd17: 256'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd18: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd19: 256'b0000000000000000000000000001011100000001000101110011111111111111000000010011111101111111111111110111111111111111111111111111111100000111011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd20: 256'b0000001101111111011111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd21: 256'b0000000000000000000000000000000100000000000000110001011101111111000000000001011100010111111111110001111111111111111111111111111100000001000111110011111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd22: 256'b0000000000000000000000000000000000000000000000010000000100011111000000000000000100000011011111110001011101111111011111111111111100000000000001110001011101111111000101111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111;
		6'd23: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000101110000000000000001000000010001011100000001001111110111111111111111;
		6'd24: 256'b0000000100010111000101111111111100111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd25: 256'b0000000000000000000000000000000000000000000000010000000100010111000000000000000100000001001111110000011101111111011111111111111100000000000000110001011101111111000101110111111111111111111111110001111111111111111111111111111111111111111111111111111111111111;
		6'd26: 256'b0000000000000000000000000000000000000000000000000000000000000111000000000000000000000001000101110000000100010111001111111111111100000000000000010000000100011111000000110111111101111111111111110001011101111111011111111111111111111111111111111111111111111111;
		6'd27: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000101110001011101111111;
		6'd28: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000111000101110111111100000000000000000000000000000111000000010001011100010111111111110000000100011111001111111111111101111111111111111111111111111111;
		6'd29: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000100111111;
		6'd30: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111;
		6'd31: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd32: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd33: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd34: 256'b0000011101111111011111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd35: 256'b0000000000000000000000000000000100000000000001110001011101111111000000010001011100010111111111110011111111111111111111111111111100000001001111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd36: 256'b0000000100010111000111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd37: 256'b0000000000000000000000000000000000000000000000010000000100011111000000000000000100000011011111110001011101111111011111111111111100000000000001110001011101111111000101111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111;
		6'd38: 256'b0000000000000000000000000000000000000000000000000000000000010111000000000000000000000001000101110000000100011111011111111111111100000000000000010000000100111111000001110111111101111111111111110001011101111111111111111111111111111111111111111111111111111111;
		6'd39: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011100000000000101110001011111111111;
		6'd40: 256'b0000000000000001000001110111111100010111011111110111111111111111000101111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd41: 256'b0000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000101110000000100010111000111111111111100000000000000010000000100010111000000010111111101111111111111110000011101111111011111111111111111111111111111111111111111111111;
		6'd42: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000011000101110111111100000000000000000000000000000111000000010001011100010111111111110000000100011111001111111111111101111111111111111111111111111111;
		6'd43: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000100111111;
		6'd44: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001011100000000000000000000000000000001000000000000000100000011011111110000000000000111000101110111111100010111111111111111111111111111;
		6'd45: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111;
		6'd46: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd47: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd48: 256'b0000000000000000000000000001011100000001000101110001111111111111000000010011111101111111111111110111111111111111111111111111111100000111011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd49: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000110111111100000000000000000000000000000001000000000000011100010111011111110000000100010111000101111111111100111111111111111111111111111111;
		6'd50: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001011100000000000000000000000000000001000000000000000100000001001111110000000000000001000001110111111100010111011111111111111111111111;
		6'd51: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
		6'd52: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000101110000000000000000000000010001011100000001001111110111111111111111;
		6'd53: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd54: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd55: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd56: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000101110001011101111111;
		6'd57: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd58: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd59: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd60: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd61: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd62: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd63: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return msg_bit_ind;
endfunction

function SubcodeInstruction page_1_get_instruction(UInt#(6) instr_counter);
	SubcodeInstruction ci;
	ci.offset = 0;
	ci.instructionVector = replicate(R1N256);
	case (instr_counter)
		6'd0 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd1 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd2 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd3 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd4 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd5 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd6 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd7 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = ML2N16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; end
		6'd8 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd9 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd10 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd11 : begin ci.offset = 28; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = R1N16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = REPR04N8; ci.instructionVector[10] = SPCN16; end
		6'd12 : begin ci.offset = 62; ci.instructionVector[0] = R14SPCN8; end
		6'd13 : begin ci.offset = 28; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = R1N32; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPR04N8; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = ML2N8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = SPCN16; end
		6'd14 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = ML2R04N8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = ML2N16; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = R0N16; end
		6'd15 : begin ci.offset = 6; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = ML2R04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = ML2N8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = R0N64; end
		6'd16 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd17 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd18 : begin ci.offset = 62; ci.instructionVector[0] = R14SPCN8; end
		6'd19 : begin ci.offset = 28; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = R14SPCN8; ci.instructionVector[9] = SPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = R0N16; end
		6'd20 : begin ci.offset = 56; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; end
		6'd21 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = ML2N8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPR04N8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N16; end
		6'd22 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = R1N8; ci.instructionVector[3] = R14SPCN8; ci.instructionVector[4] = R1N8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = R1N16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPR04N8; ci.instructionVector[13] = ML2R04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = ML2N8; ci.instructionVector[16] = SPCN8; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N16; end
		6'd23 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = ML2R04N8; ci.instructionVector[3] = R14SPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPR04N8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd24 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; end
		6'd25 : begin ci.offset = 12; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = R1N8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = ML2R04N8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = R14SPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N32; end
		6'd26 : begin ci.offset = 12; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = ML2N8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = R0N16; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = R0N32; end
		6'd27 : begin ci.offset = 2; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = R0N8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = R0N32; ci.instructionVector[12] = R0N64; end
		6'd28 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = ML2N8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = R1N8; ci.instructionVector[5] = R14SPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = R0N8; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd29 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = ML2R04N8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = R0N64; ci.instructionVector[6] = R0N128; end
		6'd30 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd31 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd32 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd33 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd34 : begin ci.offset = 52; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = ML2R04N8; end
		6'd35 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = ML2N16; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = R1N8; ci.instructionVector[8] = R14SPCN8; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = R0N8; ci.instructionVector[13] = REPN8; ci.instructionVector[14] = REPR04N8; ci.instructionVector[15] = ML2R04N8; ci.instructionVector[16] = R0N8; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; end
		6'd36 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = ML2N16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; end
		6'd37 : begin ci.offset = 14; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = R1N8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPR04N8; ci.instructionVector[11] = ML2N8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N32; end
		6'd38 : begin ci.offset = 8; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = ML2R04N8; ci.instructionVector[6] = R14SPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = ML2N16; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = R0N16; ci.instructionVector[15] = REPR04N8; ci.instructionVector[16] = R0N8; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = R0N32; end
		6'd39 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = R0N32; ci.instructionVector[12] = R0N64; end
		6'd40 : begin ci.offset = 30; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = SPCN8; ci.instructionVector[10] = SPCN16; end
		6'd41 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = ML2R04N8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = R14SPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = R1N8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = REPR04N8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd42 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = R14SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = ML2R04N8; ci.instructionVector[10] = R0N8; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = ML2R04N8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd43 : begin ci.offset = 0; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd44 : begin ci.offset = 4; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = ML2N8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd45 : begin ci.offset = 0; ci.instructionVector[0] = REPR04N8; ci.instructionVector[1] = R0N8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd46 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd47 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd48 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = ML2N16; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = R0N8; ci.instructionVector[13] = ML2R04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = R0N16; end
		6'd49 : begin ci.offset = 6; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = R14SPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = SPCN16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd50 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = ML2N8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd51 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd52 : begin ci.offset = 2; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd53 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd54 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd55 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd56 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = ML2R04N8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = R0N128; end
		6'd57 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd58 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd59 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd60 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd61 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd62 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd63 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
	endcase
	return ci;
endfunction

function Codeword page_1_get_msg_bit_ind(UInt#(6) subcodeword_counter);
	Codeword msg_bit_ind=case (subcodeword_counter)
		6'd0: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd3: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd4: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd5: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd6: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd7: 256'b0000000100010111000101111111111100111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd8: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd9: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd10: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd11: 256'b0000000000000001000001110111111100010111011111111111111111111111000101111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd12: 256'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd13: 256'b0000000000000001000000010001011100000001001111110111111111111111000001110111111101111111111111111111111111111111111111111111111100010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd14: 256'b0000000000000000000000000000011100000001000101110001011111111111000000010001111100111111111111110111111111111111111111111111111100000011011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd15: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000010011111100000000000000000000000000000001000000000000001100000111011111110000000000010111000101110111111100011111111111111111111111111111;
		6'd16: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd17: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd18: 256'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd19: 256'b0000000000000000000000010001011100000001000111110111111111111111000000110111111101111111111111110111111111111111111111111111111100010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd20: 256'b0000011101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd21: 256'b0000000000000000000000000000000100000000000001110001011101111111000000010001011100011111111111110111111111111111111111111111111100000001001111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd22: 256'b0000000000000000000000000000000100000000000000010000000100111111000000000000001100000111011111110001011101111111111111111111111100000000000101110001011111111111000111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd23: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001000101110000000000000001000000010001111100000011011111110111111111111111;
		6'd24: 256'b0000000100010111000111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd25: 256'b0000000000000000000000000000000000000000000000010000000100011111000000000000000100000011011111110001011101111111011111111111111100000000000001110001011101111111000101111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111;
		6'd26: 256'b0000000000000000000000000000000000000000000000000000000000010111000000000000000000000001000101110000000100011111011111111111111100000000000000010000000100111111000001110111111101111111111111110001011101111111111111111111111111111111111111111111111111111111;
		6'd27: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011100000000000101110001011111111111;
		6'd28: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000111000101110111111100000000000000000000000000010111000000010001011100011111111111110000000100111111011111111111111101111111111111111111111111111111;
		6'd29: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000001101111111;
		6'd30: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111;
		6'd31: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd32: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd33: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd34: 256'b0000001101111111011111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd35: 256'b0000000000000000000000000000000100000000000000110000011101111111000000000001011100010111111111110001111111111111111111111111111100000001000111110011111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd36: 256'b0000000100010111000111111111111100111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd37: 256'b0000000000000000000000000000000000000000000000010000000100010111000000000000000100000001001111110000011101111111011111111111111100000000000000110001011101111111000101111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111;
		6'd38: 256'b0000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000101110000000100010111001111111111111100000000000000010000000100011111000000110111111101111111111111110001011101111111011111111111111111111111111111111111111111111111;
		6'd39: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000001110001011101111111;
		6'd40: 256'b0000000000000001000000010111111100000111011111110111111111111111000101110111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd41: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001110000000000010111000101111111111100000000000000000000000100010111000000010001111101111111111111110000001101111111011111111111111101111111111111111111111111111111;
		6'd42: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000001000000110111111100000000000000000000000000000011000000000000011100010111011111110000000100010111000111111111111101111111111111111111111111111111;
		6'd43: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100011111;
		6'd44: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001011100000000000000000000000000000001000000000000000100000001001111110000000000000001000001110111111100010111011111111111111111111111;
		6'd45: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
		6'd46: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd47: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd48: 256'b0000000000000000000000000000001100000000000101110001011111111111000000010001011100111111111111110111111111111111111111111111111100000001011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd49: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001111100000000000000000000000000000001000000000000000100000111011111110000000000000111000101110111111100010111111111111111111111111111;
		6'd50: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000100000001000101110000000000000001000000010011111100000111011111110111111111111111;
		6'd51: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd52: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000110000000000000000000000000001011100000001000101110001111111111111;
		6'd53: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd54: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd55: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd56: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000110001011101111111;
		6'd57: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd58: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd59: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd60: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd61: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd62: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd63: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return msg_bit_ind;
endfunction

function SubcodeInstruction page_2_get_instruction(UInt#(6) instr_counter);
	SubcodeInstruction ci;
	ci.offset = 0;
	ci.instructionVector = replicate(R1N256);
	case (instr_counter)
		6'd0 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd1 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd2 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd3 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd4 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd5 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd6 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd7 : begin ci.offset = 44; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = ML2N16; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = SPCN8; end
		6'd8 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd9 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd10 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd11 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = ML2N16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = R1N8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPR04N8; ci.instructionVector[10] = R0N8; end
		6'd12 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd13 : begin ci.offset = 30; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = ML2N8; ci.instructionVector[9] = SPCN8; ci.instructionVector[10] = SPCN16; end
		6'd14 : begin ci.offset = 24; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R1N16; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = ML2N8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = ML2N16; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = R0N8; ci.instructionVector[13] = R0N16; end
		6'd15 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = R14SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = ML2R04N8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = R0N32; end
		6'd16 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd17 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd18 : begin ci.offset = 60; ci.instructionVector[0] = ML2N16; end
		6'd19 : begin ci.offset = 30; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = ML2N8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; ci.instructionVector[10] = SPCN16; end
		6'd20 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd21 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = ML2N16; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = R0N8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = R0N16; end
		6'd22 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = ML2N16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = R1N16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPR04N8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = ML2R04N8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; end
		6'd23 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = ML2N8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd24 : begin ci.offset = 44; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = ML2N16; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = SPCN8; end
		6'd25 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = R1N8; ci.instructionVector[3] = R14SPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = R1N16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = ML2R04N8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = R14SPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; end
		6'd26 : begin ci.offset = 12; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = ML2N8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = R0N16; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = R0N32; end
		6'd27 : begin ci.offset = 2; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = R0N32; ci.instructionVector[12] = R0N64; end
		6'd28 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = ML2N8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = R1N8; ci.instructionVector[5] = R14SPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = R0N8; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd29 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = ML2R04N8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = R0N32; ci.instructionVector[8] = R0N128; end
		6'd30 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd31 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd32 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd33 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd34 : begin ci.offset = 52; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = ML2R04N8; end
		6'd35 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = R1N16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPR04N8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPR04N8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; end
		6'd36 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = ML2N16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = R0N8; end
		6'd37 : begin ci.offset = 14; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPR04N8; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = ML2R04N8; ci.instructionVector[10] = R14SPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = SPCN16; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = R0N32; end
		6'd38 : begin ci.offset = 8; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = ML2N8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R1N8; ci.instructionVector[10] = R14SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = ML2R04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd39 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = ML2R04N8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = R0N32; ci.instructionVector[12] = R0N64; end
		6'd40 : begin ci.offset = 30; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = ML2R04N8; ci.instructionVector[8] = R14SPCN8; ci.instructionVector[9] = SPCN8; ci.instructionVector[10] = SPCN16; end
		6'd41 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = ML2N8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = R1N8; ci.instructionVector[5] = R14SPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = R0N8; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = R0N8; ci.instructionVector[15] = ML2R04N8; ci.instructionVector[16] = R0N8; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd42 : begin ci.offset = 6; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = ML2R04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = ML2N8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = R0N64; end
		6'd43 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd44 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = R14SPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd45 : begin ci.offset = 0; ci.instructionVector[0] = ML2R04N8; ci.instructionVector[1] = R0N8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd46 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd47 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd48 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = ML2N16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPR04N8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N16; end
		6'd49 : begin ci.offset = 4; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = ML2N8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = SPCN16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd50 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = ML2N8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = R14SPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPR04N8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd51 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd52 : begin ci.offset = 2; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPR04N8; ci.instructionVector[4] = R0N8; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = R0N32; ci.instructionVector[12] = R0N64; end
		6'd53 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd54 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd55 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd56 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = ML2R04N8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = R0N32; ci.instructionVector[8] = R0N128; end
		6'd57 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd58 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd59 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd60 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd61 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd62 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd63 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
	endcase
	return ci;
endfunction

function Codeword page_2_get_msg_bit_ind(UInt#(6) subcodeword_counter);
	Codeword msg_bit_ind=case (subcodeword_counter)
		6'd0: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd3: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd4: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd5: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd6: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd7: 256'b0000000100011111001111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd8: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd9: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd10: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd11: 256'b0000000000000111000101110111111100010111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd12: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd13: 256'b0000000000000001000000010011111100000111011111110111111111111111000101110111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd14: 256'b0000000000000000000000000001011100000001000101110011111111111111000000010011111101111111111111110111111111111111111111111111111100010111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd15: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000001000000110111111100000000000000000000000000000001000000000000011100010111011111110000000100010111000111111111111101111111111111111111111111111111;
		6'd16: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd17: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd18: 256'b0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd19: 256'b0000000000000001000000010001011100000001001111110111111111111111000001110111111101111111111111111111111111111111111111111111111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd20: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd21: 256'b0000000000000000000000000000011100000000000101110001011111111111000000010001011100111111111111110111111111111111111111111111111100000001011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd22: 256'b0000000000000000000000000000000100000000000000010000001101111111000000000000011100010111011111110001011111111111111111111111111100000001000101110001111111111111001111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd23: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000100000001000101110000000000000001000000010011111100000111011111110111111111111111;
		6'd24: 256'b0000000100010111001111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd25: 256'b0000000000000000000000000000000100000000000000010000000100011111000000000000000100000011011111110001011101111111111111111111111100000000000101110001011101111111000111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd26: 256'b0000000000000000000000000000000000000000000000000000000000010111000000000000000000000001000101110000000100011111011111111111111100000000000000010000000100111111000001110111111101111111111111110001011101111111111111111111111111111111111111111111111111111111;
		6'd27: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011100000001000101110001011111111111;
		6'd28: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000111000101110111111100000000000000000000000000010111000000010001011100011111111111110000000100111111011111111111111101111111111111111111111111111111;
		6'd29: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010000001101111111;
		6'd30: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010111;
		6'd31: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd32: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd33: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd34: 256'b0000001101111111011111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd35: 256'b0000000000000000000000000000000100000000000000010000011101111111000000000000011100010111011111110001011111111111111111111111111100000001000101110001111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd36: 256'b0000000000010111000101111111111100111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd37: 256'b0000000000000000000000000000000000000000000000000000000100010111000000000000000100000001000111110000001101111111011111111111111100000000000000010000011101111111000101110111111111111111111111110001111111111111111111111111111111111111111111111111111111111111;
		6'd38: 256'b0000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000101110000000100010111000111111111111100000000000000010000000100010111000000010011111101111111111111110000011101111111011111111111111111111111111111111111111111111111;
		6'd39: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000110001011101111111;
		6'd40: 256'b0000000000000001000000010001111100000011011111110111111111111111000101110111111111111111111111111111111111111111111111111111111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd41: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000110000000000010111000101110111111100000000000000000000000000010111000000010001011100011111111111110000000100111111011111111111111101111111111111111111111111111111;
		6'd42: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000010011111100000000000000000000000000000001000000000000001100010111011111110000000000010111000101111111111100011111111111111111111111111111;
		6'd43: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010111;
		6'd44: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001011100000000000000000000000000000000000000000000000100000001000111110000000000000001000000010111111100000111011111110111111111111111;
		6'd45: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
		6'd46: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd47: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd48: 256'b0000000000000000000000000000000100000000000001110001011101111111000000010001011100010111111111110011111111111111111111111111111100000001000111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd49: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001011100000000000000000000000000000001000000000000000100000001001111110000000000000001000001110111111100010111011111111111111111111111;
		6'd50: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001000101110000000000000001000000010001111100000001001111110111111111111111;
		6'd51: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd52: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011100000001000101110001011111111111;
		6'd53: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd54: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd55: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd56: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010000001101111111;
		6'd57: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd58: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd59: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd60: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd61: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd62: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd63: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return msg_bit_ind;
endfunction

function SubcodeInstruction page_3_get_instruction(UInt#(6) instr_counter);
	SubcodeInstruction ci;
	ci.offset = 0;
	ci.instructionVector = replicate(R1N256);
	case (instr_counter)
		6'd0 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd1 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd2 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd3 : begin ci.offset = 62; ci.instructionVector[0] = R14SPCN8; end
		6'd4 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd5 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd6 : begin ci.offset = 52; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; end
		6'd7 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPR04N8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = ML2N8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = R1N8; ci.instructionVector[12] = R14SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = SPCN8; ci.instructionVector[17] = R0N16; end
		6'd8 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd9 : begin ci.offset = 44; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; end
		6'd10 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = SPCN8; end
		6'd11 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = R1N16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = ML2R04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N16; end
		6'd12 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = R1N8; ci.instructionVector[6] = R14SPCN8; ci.instructionVector[7] = R1N8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; end
		6'd13 : begin ci.offset = 14; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = ML2R04N8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N32; end
		6'd14 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = ML2N16; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = REPR04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd15 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = ML2R04N8; ci.instructionVector[5] = R0N8; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd16 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd17 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = ML2N16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; end
		6'd18 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = R1N16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = R0N8; end
		6'd19 : begin ci.offset = 8; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = ML2R04N8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = REPN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = SPCN8; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = R0N32; end
		6'd20 : begin ci.offset = 28; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = ML2R04N8; ci.instructionVector[10] = ML2N8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = SPCN16; end
		6'd21 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = ML2N16; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = REPR04N8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd22 : begin ci.offset = 6; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = R0N64; end
		6'd23 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd24 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = ML2N8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = ML2R04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = R0N16; end
		6'd25 : begin ci.offset = 4; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = R0N8; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = ML2R04N8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = R0N32; ci.instructionVector[15] = R0N64; end
		6'd26 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = ML2R04N8; ci.instructionVector[3] = R14SPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPR04N8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd27 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd28 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = R0N8; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd29 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd30 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd31 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd32 : begin ci.offset = 62; ci.instructionVector[0] = REPSPCN8; end
		6'd33 : begin ci.offset = 24; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R1N16; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = ML2R04N8; ci.instructionVector[11] = R14SPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; end
		6'd34 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPR04N8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = ML2N8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = R1N8; ci.instructionVector[12] = R14SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = R0N8; ci.instructionVector[17] = R0N16; end
		6'd35 : begin ci.offset = 6; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = R0N16; ci.instructionVector[16] = R0N64; end
		6'd36 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = ML2N16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = R1N16; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = R0N8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPR04N8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; end
		6'd37 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd38 : begin ci.offset = 2; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd39 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd40 : begin ci.offset = 8; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPR04N8; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = REPN16; ci.instructionVector[10] = R14SPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = R0N8; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = R0N32; end
		6'd41 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = R0N8; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd42 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = ML2R04N8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = R0N64; ci.instructionVector[6] = R0N128; end
		6'd43 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd44 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd45 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd46 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd47 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd48 : begin ci.offset = 4; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = R14SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = ML2R04N8; ci.instructionVector[10] = R0N8; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = R0N64; end
		6'd49 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd50 : begin ci.offset = 0; ci.instructionVector[0] = REPR04N8; ci.instructionVector[1] = R0N8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd51 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd52 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd53 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd54 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd55 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd56 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd57 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd58 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd59 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd60 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd61 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd62 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd63 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
	endcase
	return ci;
endfunction

function Codeword page_3_get_msg_bit_ind(UInt#(6) subcodeword_counter);
	Codeword msg_bit_ind=case (subcodeword_counter)
		6'd0: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd3: 256'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd4: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd5: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd6: 256'b0001011101111111011111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd7: 256'b0000000000000000000000010001011100000001000101110001111111111111000000010011111101111111111111110111111111111111111111111111111100000111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd8: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd9: 256'b0001011101111111011111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd10: 256'b0000000101111111011111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd11: 256'b0000000000000000000000000000000100000000000000110001011101111111000000000001011100010111011111110001011111111111111111111111111100000001000101110001111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd12: 256'b0000000100010111000101111111111100011111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd13: 256'b0000000000000000000000000000000000000000000000010000000100010111000000000000000100000011011111110001011101111111011111111111111100000000000001110001011101111111000101110111111101111111111111110001011111111111111111111111111111111111111111111111111111111111;
		6'd14: 256'b0000000000000000000000000000000000000000000000000000000000000111000000000000000000000001000101110000000100010111001111111111111100000000000000010000000100011111000000110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd15: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001100000000000101110001011101111111;
		6'd16: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd17: 256'b0000000100010111000111111111111100111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd18: 256'b0000000000010111000101110111111100010111011111111111111111111111000111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd19: 256'b0000000000000000000000000000000000000000000000000000000100010111000000000000000100000001000101110000000101111111011111111111111100000000000000010000001101111111000101110111111101111111111111110001011101111111011111111111111111111111111111111111111111111111;
		6'd20: 256'b0000000000000001000000010011111100000011011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd21: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001110000000000010111000101110111111100000000000000000000000100010111000000010001011100111111111111110000000101111111011111111111111101111111111111111111111111111111;
		6'd22: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000010111111100000000000000000000000000000001000000000000011100010111011111110000000100010111000101110111111100011111111111111111111111111111;
		6'd23: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111;
		6'd24: 256'b0000000000000000000000000000001100000000000101110001011101111111000000010001011100011111111111110111111111111111111111111111111100000001001111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd25: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001011100000000000000000000000000000001000000000000000100000011011111110000000000000111000101110111111100010111011111111111111111111111;
		6'd26: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000001000101110000000000000001000000010001111100000011011111110111111111111111;
		6'd27: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd28: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011100000001000101110001011101111111;
		6'd29: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd30: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd31: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd32: 256'b0001011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd33: 256'b0000000000000001000000010001111100000011011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd34: 256'b0000000000000000000000000001011100000001000101110001111111111111000000010011111101111111111111110111111111111111111111111111111100000111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd35: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000010111111100000000000000000000000000000001000000000000011100010111011111110000000100010111000101110111111100011111111111111111111111111111;
		6'd36: 256'b0000000000000000000000000000000100000000000000010000011101111111000000000001011100010111011111110001011101111111111111111111111100000001000101110001011111111111001111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd37: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000100000001000101110000000000000001000000010111111100000111011111110111111111111111;
		6'd38: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001110000000000000000000000010001011100000001000101110001111111111111;
		6'd39: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd40: 256'b0000000000000000000000000000000000000000000000000000000000010111000000000000000100000001000101110000000100011111011111111111111100000000000000010000000101111111000001110111111101111111111111110001011101111111011111111111111111111111111111111111111111111111;
		6'd41: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011100000000000101110001011101111111;
		6'd42: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000001101111111;
		6'd43: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd44: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111;
		6'd45: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd46: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd47: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd48: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000001110111111100000000000000000000000000000011000000000001011100010111011111110000000100010111000111111111111100111111111111111111111111111111;
		6'd49: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010111;
		6'd50: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
		6'd51: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd52: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd53: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd54: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd55: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd56: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd57: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd58: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd59: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd60: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd61: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd62: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd63: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return msg_bit_ind;
endfunction

function SubcodeInstruction page_4_get_instruction(UInt#(6) instr_counter);
	SubcodeInstruction ci;
	ci.offset = 0;
	ci.instructionVector = replicate(R1N256);
	case (instr_counter)
		6'd0 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd1 : begin ci.offset = 62; ci.instructionVector[0] = R14SPCN8; end
		6'd2 : begin ci.offset = 60; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; end
		6'd3 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; end
		6'd4 : begin ci.offset = 44; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; end
		6'd5 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPR04N8; ci.instructionVector[17] = R0N8; end
		6'd6 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; end
		6'd7 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = ML2R04N8; ci.instructionVector[4] = ML2N16; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = REPSPCN8; ci.instructionVector[18] = R0N8; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd8 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; end
		6'd9 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPR04N8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = ML2N8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; end
		6'd10 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = R1N8; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = SPCN8; ci.instructionVector[18] = SPCN16; end
		6'd11 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = R0N8; ci.instructionVector[13] = R0N16; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = ML2R04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = SPCN16; ci.instructionVector[21] = R0N16; ci.instructionVector[22] = R0N32; end
		6'd12 : begin ci.offset = 12; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = REPN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = REPN8; ci.instructionVector[17] = REPSPCN8; ci.instructionVector[18] = REPSPCN8; ci.instructionVector[19] = R0N8; ci.instructionVector[20] = SPCN16; ci.instructionVector[21] = R0N16; end
		6'd13 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = ML2R04N8; ci.instructionVector[6] = R0N8; ci.instructionVector[7] = ML2N8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = R0N32; ci.instructionVector[16] = R0N64; end
		6'd14 : begin ci.offset = 2; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = ML2R04N8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd15 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd16 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = R1N8; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; end
		6'd17 : begin ci.offset = 14; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = REPN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = REPSPCN8; ci.instructionVector[18] = SPCN8; ci.instructionVector[19] = ML2R04N8; ci.instructionVector[20] = R0N8; ci.instructionVector[21] = R0N16; end
		6'd18 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPR04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = REPN8; ci.instructionVector[19] = SPCN8; ci.instructionVector[20] = SPCN16; ci.instructionVector[21] = SPCN16; ci.instructionVector[22] = R0N16; end
		6'd19 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = ML2R04N8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd20 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPR04N8; ci.instructionVector[7] = R14SPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R1N8; ci.instructionVector[11] = R14SPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = REPSPCN8; ci.instructionVector[18] = SPCN8; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd21 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = SPCN16; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd22 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = ML2R04N8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = R0N32; ci.instructionVector[8] = R0N128; end
		6'd23 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd24 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = R0N8; ci.instructionVector[13] = R0N16; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPR04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = SPCN16; ci.instructionVector[21] = R0N16; ci.instructionVector[22] = R0N32; end
		6'd25 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = R0N64; ci.instructionVector[6] = R0N128; end
		6'd26 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = R0N8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd27 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd28 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd29 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd30 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd31 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd32 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPR04N8; ci.instructionVector[16] = SPCN16; end
		6'd33 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = REPSPCN8; ci.instructionVector[18] = SPCN8; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd34 : begin ci.offset = 4; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = REPR04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = SPCN16; ci.instructionVector[20] = R0N16; ci.instructionVector[21] = R0N32; end
		6'd35 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = R0N32; ci.instructionVector[8] = R0N128; end
		6'd36 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R0N8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPR04N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = R0N64; end
		6'd37 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd38 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd39 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd40 : begin ci.offset = 2; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd41 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd42 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd43 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd44 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd45 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd46 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd47 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd48 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = R0N32; ci.instructionVector[8] = R0N128; end
		6'd49 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd50 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd51 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd52 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd53 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd54 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd55 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd56 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd57 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd58 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd59 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd60 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd61 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd62 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd63 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
	endcase
	return ci;
endfunction

function Codeword page_4_get_msg_bit_ind(UInt#(6) subcodeword_counter);
	Codeword msg_bit_ind=case (subcodeword_counter)
		6'd0: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1: 256'b0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2: 256'b0001011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd3: 256'b0000000100010111000101110111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd4: 256'b0001011101111111011111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd5: 256'b0000000000000111000101110111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd6: 256'b0000000000000001000000010111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd7: 256'b0000000000000000000000000000000000000000000000000000000000010111000000000000000100000001000101110000000100010111000101110111111100000000000000010000000100010111000000010001011100111111111111110000001101111111011111111111111101111111111111111111111111111111;
		6'd8: 256'b0001011101111111011111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd9: 256'b0000000000000001000000010001011100000001001111110111111111111111000001110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd10: 256'b0000000000000001000000010001011100000001000101110001011101111111000000010001011100011111111111110111111111111111111111111111111100000001011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd11: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000011000101110111111100000000000000000000000000010111000000010001011100010111011111110000000100010111000101110111111100010111011111110111111111111111;
		6'd12: 256'b0000000000000000000000000000000100000000000101110001011101111111000000010001011100010111011111110001011101111111011111111111111100000001000101110001011101111111000101110111111101111111111111110001011101111111111111111111111111111111111111111111111111111111;
		6'd13: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001011100000000000000000000000000000001000000000000000100000001001111110000000000000011000101110111111100010111011111110111111111111111;
		6'd14: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000001000101110000000000000001000000010001011100000001000101110001111111111111;
		6'd15: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd16: 256'b0000000100010111000111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd17: 256'b0000000000000000000000000000001100000001000101110001011101111111000000010001011100010111011111110001011101111111011111111111111100000001000101110001011101111111000101110111111111111111111111110001111111111111111111111111111111111111111111111111111111111111;
		6'd18: 256'b0000000000000000000000000000000100000000000000010000000101111111000000000000011100010111011111110001011101111111011111111111111100000001000101110001011101111111000101110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd19: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001011100000000000000000000000000000000000000000000000100000001000101110000000000000001000000010001011100000011011111110111111111111111;
		6'd20: 256'b0000000000000000000000000000000000000000000000000000000100010111000000000000000100000001000101110000000100010111000111111111111100000000000000010000000100011111000001110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd21: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000000000000010001011100000001000101110001011101111111;
		6'd22: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010000001101111111;
		6'd23: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd24: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000111000101110111111100000000000000000000000000010111000000010001011100010111011111110000000100010111000101110111111100010111011111110111111111111111;
		6'd25: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000100010111;
		6'd26: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111;
		6'd27: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd28: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd29: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd30: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd31: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd32: 256'b0000000000000001000001110111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd33: 256'b0000000000000000000000000000000000000000000000000000000100010111000000000000000100000001000101110000000100010111000101110111111100000000000000010000000100010111000000010111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd34: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001110000000100010111000101110111111100000000000000000000000100010111000000010001011100010111011111110000000100010111000101111111111100111111111111111111111111111111;
		6'd35: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010000000101111111;
		6'd36: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000010001011100000000000000000000000000000001000000000000000100000111011111110000000000010111000101110111111100010111011111110111111111111111;
		6'd37: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111;
		6'd38: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd39: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd40: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000101110000000000000001000000010001011100000001000101110001011111111111;
		6'd41: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd42: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd43: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd44: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd45: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd46: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd47: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd48: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010001011101111111;
		6'd49: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd50: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd51: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd52: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd53: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd54: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd55: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd56: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd57: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd58: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd59: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd60: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd61: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd62: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd63: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return msg_bit_ind;
endfunction

function SubcodeInstruction page_5_get_instruction(UInt#(6) instr_counter);
	SubcodeInstruction ci;
	ci.offset = 0;
	ci.instructionVector = replicate(R1N256);
	case (instr_counter)
		6'd0 : begin ci.offset = 0; ci.instructionVector[0] = R1N256; end
		6'd1 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd2 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd3 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = ML2N16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = R1N8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; end
		6'd4 : begin ci.offset = 60; ci.instructionVector[0] = REPN16; end
		6'd5 : begin ci.offset = 30; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = R0N8; end
		6'd6 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = SPCN16; end
		6'd7 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R1N8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = REPR04N8; ci.instructionVector[18] = R0N8; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd8 : begin ci.offset = 44; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; end
		6'd9 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = ML2N8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = SPCN16; end
		6'd10 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPR04N8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = ML2N8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = R1N8; ci.instructionVector[12] = R14SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = SPCN8; ci.instructionVector[17] = SPCN16; end
		6'd11 : begin ci.offset = 6; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = REPR04N8; ci.instructionVector[10] = R0N8; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = SPCN16; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = R0N32; end
		6'd12 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = R1N8; ci.instructionVector[3] = R14SPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = REPN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = REPR04N8; ci.instructionVector[18] = R0N8; ci.instructionVector[19] = SPCN16; ci.instructionVector[20] = R0N16; end
		6'd13 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPR04N8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = R0N16; ci.instructionVector[14] = R0N32; ci.instructionVector[15] = R0N64; end
		6'd14 : begin ci.offset = 2; ci.instructionVector[0] = R14SPCN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = R0N8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd15 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd16 : begin ci.offset = 28; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = R1N16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = ML2N8; ci.instructionVector[8] = SPCN8; end
		6'd17 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = R1N8; ci.instructionVector[4] = R14SPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = R1N16; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N16; end
		6'd18 : begin ci.offset = 12; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = REPN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = ML2R04N8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = ML2N8; ci.instructionVector[17] = SPCN8; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = SPCN16; ci.instructionVector[20] = R0N16; end
		6'd19 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = ML2N8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = R0N16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = R0N32; ci.instructionVector[13] = R0N64; end
		6'd20 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = ML2R04N8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R1N8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = REPR04N8; ci.instructionVector[18] = R0N8; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd21 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = R0N128; end
		6'd22 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = R0N64; ci.instructionVector[6] = R0N128; end
		6'd23 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd24 : begin ci.offset = 4; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = R0N8; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = SPCN16; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = R0N64; end
		6'd25 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd26 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd27 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd28 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd29 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd30 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd31 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd32 : begin ci.offset = 20; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = R1N16; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN16; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPN16; ci.instructionVector[10] = REPN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPR04N8; ci.instructionVector[14] = SPCN16; end
		6'd33 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R1N8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = R0N16; ci.instructionVector[17] = REPR04N8; ci.instructionVector[18] = R0N8; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd34 : begin ci.offset = 4; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = R0N8; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPR04N8; ci.instructionVector[15] = R0N8; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N16; ci.instructionVector[20] = R0N32; end
		6'd35 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd36 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = ML2R04N8; ci.instructionVector[6] = R0N8; ci.instructionVector[7] = ML2N8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = R0N16; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = SPCN8; ci.instructionVector[14] = R0N16; ci.instructionVector[15] = R0N32; ci.instructionVector[16] = R0N64; end
		6'd37 : begin ci.offset = 0; ci.instructionVector[0] = ML2R04N8; ci.instructionVector[1] = R0N8; ci.instructionVector[2] = R0N16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd38 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd39 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd40 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = REPR04N8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = R0N32; ci.instructionVector[11] = SPCN16; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd41 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd42 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd43 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd44 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd45 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd46 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd47 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd48 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = ML2R04N8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = R0N64; ci.instructionVector[6] = R0N128; end
		6'd49 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd50 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd51 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd52 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd53 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd54 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd55 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd56 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd57 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd58 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd59 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd60 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd61 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd62 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd63 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
	endcase
	return ci;
endfunction

function Codeword page_5_get_msg_bit_ind(UInt#(6) subcodeword_counter);
	Codeword msg_bit_ind=case (subcodeword_counter)
		6'd0: 256'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd3: 256'b0000000100010111000101110111111100010111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd4: 256'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd5: 256'b0000000000010111000101110111111100010111011111110111111111111111000101110111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd6: 256'b0000000000000001000001110111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd7: 256'b0000000000000000000000000000000000000000000000000000000000000111000000000000000000000001000101110000000100010111000101111111111100000000000000010000000100010111000000110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd8: 256'b0001011101111111011111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd9: 256'b0000000000000001000000010011111100000111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd10: 256'b0000000000000001000000010001011100000001000101110001111111111111000000010011111101111111111111110111111111111111111111111111111100000111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd11: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000001000001110111111100000000000000000000000000000111000000010001011100010111011111110000000100010111000101110111111100011111111111111111111111111111;
		6'd12: 256'b0000000000000000000000000000000100000000000001110001011101111111000000010001011100010111011111110001011101111111011111111111111100000001000101110001011101111111000111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd13: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001011100000000000000000000000000000001000000000000000100000001000101110000000000000001000001110111111100010111011111110111111111111111;
		6'd14: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000101110000000000000001000000010001011100000001000101110001111111111111;
		6'd15: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd16: 256'b0000000100111111011111111111111101111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd17: 256'b0000000000000000000000000000000100000000000101110001011101111111000000010001011100010111011111110001011101111111111111111111111100000001000101110001111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd18: 256'b0000000000000000000000000000000100000000000000010000000100111111000000000000001100010111011111110001011101111111011111111111111100000001000101110001011101111111000101110111111101111111111111110001011101111111111111111111111111111111111111111111111111111111;
		6'd19: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000101110000000000000001000000010001011100000001001111110111111111111111;
		6'd20: 256'b0000000000000000000000000000000000000000000000000000000000000111000000000000000000000001000101110000000100010111000101111111111100000000000000010000000100010111000000110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd21: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000101110001011101111111;
		6'd22: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000000100010111;
		6'd23: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd24: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000010111111100000000000000000000000000000001000000000001011100010111011111110000000100010111000101110111111100010111011111111111111111111111;
		6'd25: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010111;
		6'd26: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd27: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd28: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd29: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd30: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd31: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd32: 256'b0000000000000001000001110111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd33: 256'b0000000000000000000000000000000000000000000000000000000000000111000000000000000000000001000101110000000100010111000101111111111100000000000000010000000100010111000000010111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd34: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000111000101110111111100000000000000000000000000010111000000010001011100010111011111110000000100010111000101111111111100111111111111111111111111111111;
		6'd35: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010111;
		6'd36: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001011100000000000000000000000000000001000000000000000100000001001111110000000000000011000101110111111100010111011111110111111111111111;
		6'd37: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011;
		6'd38: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd39: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd40: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000001110000000000000000000000010001011100000001000101110001011101111111;
		6'd41: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd42: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd43: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd44: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd45: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd46: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd47: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd48: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010000001101111111;
		6'd49: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd50: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd51: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd52: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd53: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd54: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd55: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd56: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd57: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd58: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd59: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd60: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd61: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd62: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd63: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return msg_bit_ind;
endfunction

function SubcodeInstruction page_6_get_instruction(UInt#(6) instr_counter);
	SubcodeInstruction ci;
	ci.offset = 0;
	ci.instructionVector = replicate(R1N256);
	case (instr_counter)
		6'd0 : begin ci.offset = 60; ci.instructionVector[0] = ML2N16; end
		6'd1 : begin ci.offset = 30; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = R1N32; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPN16; ci.instructionVector[6] = REPN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = REPN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = SPCN8; end
		6'd2 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = SPCN8; end
		6'd3 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPR04N8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = REPN8; ci.instructionVector[19] = SPCN8; ci.instructionVector[20] = SPCN16; ci.instructionVector[21] = SPCN16; ci.instructionVector[22] = R0N16; end
		6'd4 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = REPN8; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = R0N8; end
		6'd5 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = ML2R04N8; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = REPN16; ci.instructionVector[11] = R14SPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = SPCN8; ci.instructionVector[18] = SPCN16; ci.instructionVector[19] = R0N32; end
		6'd6 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = ML2N16; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = SPCN8; ci.instructionVector[10] = SPCN16; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = SPCN8; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = REPR04N8; ci.instructionVector[19] = R0N8; ci.instructionVector[20] = R0N16; ci.instructionVector[21] = R0N32; end
		6'd7 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = R0N128; end
		6'd8 : begin ci.offset = 12; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N16; ci.instructionVector[2] = REPN16; ci.instructionVector[3] = REPN16; ci.instructionVector[4] = REPN8; ci.instructionVector[5] = REPR04N8; ci.instructionVector[6] = R1N16; ci.instructionVector[7] = REPN16; ci.instructionVector[8] = REPN16; ci.instructionVector[9] = R14SPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPN8; ci.instructionVector[12] = REPSPCN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = SPCN8; ci.instructionVector[17] = SPCN16; end
		6'd9 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = SPCN8; ci.instructionVector[18] = REPR04N8; ci.instructionVector[19] = R0N8; ci.instructionVector[20] = R0N16; ci.instructionVector[21] = SPCN16; ci.instructionVector[22] = R0N16; ci.instructionVector[23] = R0N32; end
		6'd10 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = REPN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = REPSPCN8; ci.instructionVector[6] = SPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPR04N8; ci.instructionVector[10] = R0N8; ci.instructionVector[11] = SPCN16; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = SPCN8; ci.instructionVector[15] = SPCN16; ci.instructionVector[16] = SPCN16; ci.instructionVector[17] = R0N16; ci.instructionVector[18] = R0N64; end
		6'd11 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd12 : begin ci.offset = 0; ci.instructionVector[0] = ML2N16; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = R0N32; ci.instructionVector[10] = REPSPCN8; ci.instructionVector[11] = R0N8; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd13 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd14 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd15 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd16 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN16; ci.instructionVector[2] = REPN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = REPN16; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPN8; ci.instructionVector[8] = REPSPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = REPN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPN8; ci.instructionVector[15] = REPSPCN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = R0N8; ci.instructionVector[18] = REPN8; ci.instructionVector[19] = REPSPCN8; ci.instructionVector[20] = SPCN16; ci.instructionVector[21] = SPCN16; ci.instructionVector[22] = R0N16; end
		6'd17 : begin ci.offset = 0; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = REPN8; ci.instructionVector[2] = REPR04N8; ci.instructionVector[3] = ML2N8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = SPCN8; ci.instructionVector[8] = SPCN16; ci.instructionVector[9] = SPCN16; ci.instructionVector[10] = R0N16; ci.instructionVector[11] = REPSPCN8; ci.instructionVector[12] = SPCN8; ci.instructionVector[13] = SPCN16; ci.instructionVector[14] = R0N32; ci.instructionVector[15] = R0N64; end
		6'd18 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = REPSPCN8; ci.instructionVector[3] = SPCN8; ci.instructionVector[4] = REPSPCN8; ci.instructionVector[5] = SPCN8; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = R0N8; ci.instructionVector[9] = R0N16; ci.instructionVector[10] = R0N32; ci.instructionVector[11] = SPCN16; ci.instructionVector[12] = R0N16; ci.instructionVector[13] = R0N32; ci.instructionVector[14] = R0N64; end
		6'd19 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd20 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPR04N8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = SPCN16; ci.instructionVector[4] = R0N16; ci.instructionVector[5] = SPCN16; ci.instructionVector[6] = R0N16; ci.instructionVector[7] = R0N32; ci.instructionVector[8] = R0N128; end
		6'd21 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd22 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd23 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd24 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd25 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd26 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd27 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd28 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd29 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd30 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd31 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd32 : begin ci.offset = 4; ci.instructionVector[0] = REPN16; ci.instructionVector[1] = R1N8; ci.instructionVector[2] = R14SPCN8; ci.instructionVector[3] = REPSPCN8; ci.instructionVector[4] = SPCN8; ci.instructionVector[5] = REPN8; ci.instructionVector[6] = REPSPCN8; ci.instructionVector[7] = REPSPCN8; ci.instructionVector[8] = SPCN8; ci.instructionVector[9] = REPSPCN8; ci.instructionVector[10] = SPCN8; ci.instructionVector[11] = SPCN16; ci.instructionVector[12] = REPN8; ci.instructionVector[13] = REPSPCN8; ci.instructionVector[14] = REPSPCN8; ci.instructionVector[15] = SPCN8; ci.instructionVector[16] = REPSPCN8; ci.instructionVector[17] = SPCN8; ci.instructionVector[18] = R0N16; ci.instructionVector[19] = SPCN16; ci.instructionVector[20] = R0N16; ci.instructionVector[21] = R0N32; end
		6'd33 : begin ci.offset = 0; ci.instructionVector[0] = REPN8; ci.instructionVector[1] = REPSPCN8; ci.instructionVector[2] = ML2R04N8; ci.instructionVector[3] = R0N8; ci.instructionVector[4] = SPCN16; ci.instructionVector[5] = R0N16; ci.instructionVector[6] = SPCN16; ci.instructionVector[7] = R0N16; ci.instructionVector[8] = R0N32; ci.instructionVector[9] = R0N128; end
		6'd34 : begin ci.offset = 0; ci.instructionVector[0] = REPSPCN8; ci.instructionVector[1] = SPCN8; ci.instructionVector[2] = SPCN16; ci.instructionVector[3] = R0N32; ci.instructionVector[4] = R0N64; ci.instructionVector[5] = R0N128; end
		6'd35 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd36 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd37 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd38 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd39 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd40 : begin ci.offset = 0; ci.instructionVector[0] = SPCN16; ci.instructionVector[1] = R0N16; ci.instructionVector[2] = R0N32; ci.instructionVector[3] = R0N64; ci.instructionVector[4] = R0N128; end
		6'd41 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd42 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd43 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd44 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd45 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd46 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd47 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd48 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd49 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd50 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd51 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd52 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd53 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd54 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd55 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd56 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd57 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd58 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd59 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd60 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd61 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd62 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
		6'd63 : begin ci.offset = 0; ci.instructionVector[0] = R0N256; end
	endcase
	return ci;
endfunction

function Codeword page_6_get_msg_bit_ind(UInt#(6) subcodeword_counter);
	Codeword msg_bit_ind=case (subcodeword_counter)
		6'd0: 256'b0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd1: 256'b0000000100010111000101110111111100010111011111110111111111111111000101110111111101111111111111111111111111111111111111111111111100010111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
		6'd2: 256'b0000000100010111000101110111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd3: 256'b0000000000000000000000000000000100000000000000010000000101111111000000000000011100010111011111110001011101111111011111111111111100000001000101110001011101111111000101110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd4: 256'b0000000000010111000101110111111100010111011111110111111111111111000101110111111101111111111111110111111111111111111111111111111100010111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd5: 256'b0000000000000000000000000000000000000000000000010000000100010111000000000000000100000001000101110000000100011111011111111111111100000000000000010000001101111111000101110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd6: 256'b0000000000000000000000000000000000000000000000000000000000000111000000000000000000000001000101110000000100010111000101110111111100000000000000010000000100010111000000010001011100010111011111110000000100010111001111111111111101111111111111111111111111111111;
		6'd7: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000101110001011101111111;
		6'd8: 256'b0000000000000001000000010001011100000001000101110001011101111111000000010001111101111111111111110111111111111111111111111111111100000111011111110111111111111111011111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111;
		6'd9: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001110000000100010111000101110111111100000000000000010000000100010111000000010001011100010111011111110000000100010111000101110111111100010111011111110111111111111111;
		6'd10: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000010001011100000000000000000000000000000001000000000000011100010111011111110000000100010111000101110111111100010111011111110111111111111111;
		6'd11: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010111;
		6'd12: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000100000001000101110000000000000001000000010001011100000001000101110011111111111111;
		6'd13: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd14: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd15: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd16: 256'b0000000000000000000000000000000100000000000000010001011101111111000000000001011100010111011111110001011101111111011111111111111100000001000101110001011101111111000101110111111101111111111111110001011101111111011111111111111101111111111111111111111111111111;
		6'd17: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001011100000000000000000000000000000001000000000000000100000001000101110000000000000001000000010011111100000111011111110111111111111111;
		6'd18: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000101110000000000000001000000010001011100000001000101110001011101111111;
		6'd19: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd20: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000010000011101111111;
		6'd21: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd22: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd23: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd24: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010111;
		6'd25: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd26: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd27: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd28: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd29: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd30: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd31: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd32: 256'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000101110000000100010111000101110111111100000000000000010000000100010111000000010001011100010111011111110000000100010111000111111111111101111111111111111111111111111111;
		6'd33: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000110001011101111111;
		6'd34: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100010111;
		6'd35: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd36: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd37: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd38: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd39: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd40: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		6'd41: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd42: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd43: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd44: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd45: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd46: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd47: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd48: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd49: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd50: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd51: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd52: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd53: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd54: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd55: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd56: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd57: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd58: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd59: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd60: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd61: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd62: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		6'd63: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return msg_bit_ind;
endfunction

(* noinline *)
function SubcodeInstruction get_instruction(UInt#(6) instr_counter, UInt#(3) page_num);
	SubcodeInstruction ci = case (page_num)
		3'd0: page_0_get_instruction(instr_counter);
		3'd1: page_1_get_instruction(instr_counter);
		3'd2: page_2_get_instruction(instr_counter);
		3'd3: page_3_get_instruction(instr_counter);
		3'd4: page_4_get_instruction(instr_counter);
		3'd5: page_5_get_instruction(instr_counter);
		3'd6: page_6_get_instruction(instr_counter);
	endcase;
	return ci;
endfunction

(* noinline *)
function Codeword get_msg_bit_ind(UInt#(6) subcodeword_counter, UInt#(3) page_num);
	Codeword msg_bit_ind = case (page_num)
		3'd0: page_0_get_msg_bit_ind(subcodeword_counter);
		3'd1: page_1_get_msg_bit_ind(subcodeword_counter);
		3'd2: page_2_get_msg_bit_ind(subcodeword_counter);
		3'd3: page_3_get_msg_bit_ind(subcodeword_counter);
		3'd4: page_4_get_msg_bit_ind(subcodeword_counter);
		3'd5: page_5_get_msg_bit_ind(subcodeword_counter);
		3'd6: page_6_get_msg_bit_ind(subcodeword_counter);
	endcase;
	return msg_bit_ind;
endfunction

function UInt#(6) get_msg_bit_len(UInt#(3) page_num);
	return case (page_num)
		3'd0: 6'd32;
		3'd1: 6'd32;
		3'd2: 6'd32;
		3'd3: 6'd24;
		3'd4: 6'd16;
		3'd5: 6'd16;
		3'd6: 6'd8;
	endcase;
endfunction

function UInt#(6) get_eom_bit_idx(UInt#(3) page_num);
	return case (page_num)
		3'd0: 6'd63;
		3'd1: 6'd63;
		3'd2: 6'd63;
		3'd3: 6'd63;
		3'd4: 6'd63;
		3'd5: 6'd63;
		3'd6: 6'd63;
	endcase;
endfunction
