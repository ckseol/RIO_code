function Bit#(32) get_msg_bit(UInt#(8) counter, UInt#(3) page_num);
	Bit#(32) msg_bit = case (page_num)
		3'd0: get_msg_bit_page0(truncate(counter));
		3'd1: get_msg_bit_page1(truncate(counter));
		3'd2: get_msg_bit_page2(truncate(counter));
		3'd3: get_msg_bit_page3(truncate(counter));
		3'd4: get_msg_bit_page4(truncate(counter));
		3'd5: get_msg_bit_page5(truncate(counter));
		3'd6: get_msg_bit_page6(truncate(counter));
	endcase;
	return msg_bit;
endfunction

function Bit#(32) get_msg_bit_page0(UInt#(8) counter);
	Bit#(32) out = case(counter)
		8'd0: 32'b10111011001111011110110111100100;
		8'd1: 32'b00110011111010001101100010101110;
		8'd2: 32'b01011011011110011100101011101010;
		8'd3: 32'b10001010101101001101101001111100;
		8'd4: 32'b10001000101111110110110110000100;
		8'd5: 32'b10111110011010001100011011001001;
		8'd6: 32'b01110110000110011101101100001010;
		8'd7: 32'b11111011000000011011111000111000;
		8'd8: 32'b10000010011110100111010010010010;
		8'd9: 32'b00000011110001110001010111001111;
		8'd10: 32'b10100000001100001011111000111101;
		8'd11: 32'b11111100011110010000010100000111;
		8'd12: 32'b11101001110001110000001001000011;
		8'd13: 32'b11111110010011111000100111110011;
		8'd14: 32'b00010001100101000110011101110000;
		8'd15: 32'b00000000000111001101011010101101;
		8'd16: 32'b10011001010001001110000101000010;
		8'd17: 32'b10110101111110101001101111000111;
		8'd18: 32'b00000001100111100111101000011111;
		8'd19: 32'b10100110000110110001010010111100;
		8'd20: 32'b01100100001011010011010110011110;
		8'd21: 32'b11010110110001111010001101110010;
		8'd22: 32'b00101010000100101111010110000010;
		8'd23: 32'b11101011000001001101010001010110;
		8'd24: 32'b00011011011101011111110010111000;
		8'd25: 32'b00111100010100000100110000011001;
		8'd26: 32'b01000101100110110000000000010111;
		8'd27: 32'b01100010100000111111100011010110;
		8'd28: 32'b11011100101011111000011011110011;
		8'd29: 32'b10100100100100111101011110001010;
		8'd30: 32'b11101100000001111010100101011100;
		8'd31: 32'b11100000100010011001110111011111;
		8'd32: 32'b11000111100110010101101111011001;
		8'd33: 32'b10110100100001111101101001011100;
		8'd34: 32'b11001100100111011000111000100001;
		8'd35: 32'b00001101100010101111101110111010;
		8'd36: 32'b11111111111101111100111111000101;
		8'd37: 32'b00010001001111101100011011011101;
		8'd38: 32'b01111100001110000001010100011011;
		8'd39: 32'b00010001011000110100000100100111;
		8'd40: 32'b00111100111001001000001001110101;
		8'd41: 32'b11110111011000010000001110011001;
		8'd42: 32'b10101001001111011110101110011011;
		8'd43: 32'b01011101010001111011111011010010;
		8'd44: 32'b10000000000111001110000101001110;
		8'd45: 32'b01011111011100100101110000100101;
		8'd46: 32'b10111100010111100100011100011011;
		8'd47: 32'b01010001010011001000101110000011;
		8'd48: 32'b11100100100101110001001001111000;
		8'd49: 32'b00000000011100101111100000101101;
		8'd50: 32'b01100111001000111011100011111010;
		8'd51: 32'b00010100001111010000110101101101;
		8'd52: 32'b01110100010010010010000010000010;
		8'd53: 32'b10011110111111001001110111010011;
		8'd54: 32'b00000000100000011011110000100100;
		8'd55: 32'b11100101101010000100111001010101;
		8'd56: 32'b00110111110100110100011001101001;
		8'd57: 32'b00001110001001110100111000100010;
		8'd58: 32'b01111110100010000000011100111001;
		8'd59: 32'b01100110000110001000000101001111;
		8'd60: 32'b11101000010011001100011111110001;
		8'd61: 32'b10101100100101110001100010111100;
		8'd62: 32'b00110011010111101101110000001111;
		8'd63: 32'b10100000000010011001001100101000;
		8'd64: 32'b00111110000011100101011101000011;
		8'd65: 32'b10110001110010010011000111100101;
		8'd66: 32'b01111101001111001111011001111110;
		8'd67: 32'b10100000011100010100000010111110;
		8'd68: 32'b10100101101110100111111000010101;
		8'd69: 32'b00001101001101110101110100111110;
		8'd70: 32'b01101110101010101011111111101110;
		8'd71: 32'b10000110110011100011110000111001;
		8'd72: 32'b01101000011011110100001011010010;
		8'd73: 32'b10001101010100011101010110111110;
		8'd74: 32'b01111100001110110100000101100100;
		8'd75: 32'b10010011101000000111101101010110;
		8'd76: 32'b11100100111000011110010001011100;
		8'd77: 32'b10000001010000001001101111000101;
		8'd78: 32'b10000000111110000010001000101011;
		8'd79: 32'b10010110010110110010110101100000;
		8'd80: 32'b01001001100101111000011011010100;
		8'd81: 32'b01001010010001100100001010111000;
		8'd82: 32'b10111011110010101001100110111010;
		8'd83: 32'b10101000011001011011110010011111;
		8'd84: 32'b10010111001111001000001111111011;
		8'd85: 32'b01111000111101100110011100100001;
		8'd86: 32'b00010101001000100010001111001110;
		8'd87: 32'b11111110011011111011011000011101;
		8'd88: 32'b10100100101101101000110100010101;
		8'd89: 32'b00001101010011100001101101100000;
		8'd90: 32'b01100011011001011100010010010110;
		8'd91: 32'b00011010110010000110011001100011;
		8'd92: 32'b00101111101010011110100111111000;
		8'd93: 32'b01100110110010000011001111101011;
		8'd94: 32'b01111010101110001000111100000001;
		8'd95: 32'b01110010010010111011111101011110;
		8'd96: 32'b10110101100011010110000101001001;
		8'd97: 32'b10000100010011011110001000100101;
		8'd98: 32'b01101011111001101100100100010111;
		8'd99: 32'b11010101101010110000110110111001;
		8'd100: 32'b11001001111100001000011111101100;
		8'd101: 32'b11011110111111101100000001010100;
		8'd102: 32'b10010000001011011010100000011010;
		8'd103: 32'b10011011100110111001011110101011;
		8'd104: 32'b00101111011110110101010010000010;
		8'd105: 32'b10111010110101011011111101001001;
		8'd106: 32'b00000001110000000111100001101010;
		8'd107: 32'b11010100010001110111110100001001;
		8'd108: 32'b00011000100000111101101001011111;
		8'd109: 32'b01101010111101000110001010100000;
		8'd110: 32'b11110100001100001100010001010010;
		8'd111: 32'b11000100001010101010010001001100;
		8'd112: 32'b00100100100010010000001100111101;
		8'd113: 32'b10100100000011100111000101101101;
		8'd114: 32'b10100011001001001101111000101100;
		8'd115: 32'b00011011010011101000011110110110;
		8'd116: 32'b00111111011010101101111110101101;
		8'd117: 32'b00010001111000010011101000010011;
		8'd118: 32'b11111000110111111000111000100101;
		8'd119: 32'b11101011101111100111011100110100;
		8'd120: 32'b10110000000000001000010101111100;
		8'd121: 32'b10100000001001101110001100101101;
		8'd122: 32'b10010010001011100111001010010110;
		8'd123: 32'b00101011110101110110101101000001;
		8'd124: 32'b01111001010000111010111101111000;
		8'd125: 32'b11001010010000101011111110011001;
		8'd126: 32'b11001100100111110011011011011100;
		8'd127: 32'b00101100010100110110001110101110;
		8'd128: 32'b01100011000011101001010000001011;
		8'd129: 32'b01001010100111000011100111101001;
		8'd130: 32'b11101001001101001110101101001011;
		8'd131: 32'b11010111101010010110110101100101;
		8'd132: 32'b10000000101110110100100100101101;
		8'd133: 32'b01000110010010011001001101000000;
		8'd134: 32'b11110001000000101010010000111100;
		8'd135: 32'b10001001101010110111110100001000;
		8'd136: 32'b10111001111001100100000100000100;
		8'd137: 32'b10100101111100110011001011011111;
		8'd138: 32'b11001111111100111101110101000011;
		8'd139: 32'b10001111001010000011111100010101;
		8'd140: 32'b00111000001101101101000011000101;
		8'd141: 32'b10111010101000110100000110000111;
		8'd142: 32'b01001000011111111010001101011110;
		8'd143: 32'b10011000110010000011100010001111;
		8'd144: 32'b11010010010101011100111101101101;
		8'd145: 32'b00110000110001000111001000001100;
		8'd146: 32'b01101011001100000100110000000111;
		8'd147: 32'b00110110001110110110010101110011;
		8'd148: 32'b10001001010111111011001101110110;
		8'd149: 32'b10110010111101001101010000010111;
		8'd150: 32'b11010101101101111001111001111101;
		8'd151: 32'b00100001110101011010111010100100;
		8'd152: 32'b00110111101110111011100100001100;
		8'd153: 32'b00011010101001000011100110010001;
		8'd154: 32'b00010001011000001100010100111001;
		8'd155: 32'b10010011000100100101100101111010;
		8'd156: 32'b01110111100111101101000010111000;
		8'd157: 32'b01001111001001000011111110010010;
		8'd158: 32'b11001010010101111110000011101010;
		8'd159: 32'b01101000000110001011000001101010;
		8'd160: 32'b00011011011011101001011011001100;
		8'd161: 32'b00011011101101001001100001001100;
		8'd162: 32'b10000110110011011111111010100100;
		8'd163: 32'b01100100110101110110100011001110;
		8'd164: 32'b11010111011001111011011111110101;
		8'd165: 32'b11011111111110010011000101000110;
		8'd166: 32'b01111100010001111000001000001010;
		8'd167: 32'b01001000010011101111111001000110;
		8'd168: 32'b00000111101110110101010111011000;
		8'd169: 32'b10100010101111011011011010001110;
		8'd170: 32'b11100001000001001110111010100101;
		8'd171: 32'b11110011100101010010111110111000;
		8'd172: 32'b00110011100001110000011000111010;
		8'd173: 32'b10111100110111001110110111000010;
		8'd174: 32'b10100100010101110001110000010111;
		8'd175: 32'b11001011010010110111011001110011;
		8'd176: 32'b00010010000010010001101100111100;
		8'd177: 32'b00001010001111101011010110101111;
		8'd178: 32'b10111100010110111111000000101100;
		8'd179: 32'b00110111010000100011111100011010;
		8'd180: 32'b11000010011101110101110100011111;
		8'd181: 32'b11100110110101110100110101010110;
		8'd182: 32'b01100001110001100001100010110100;
		8'd183: 32'b01011001101100000101010100011110;
		8'd184: 32'b10001101010100100000110110101111;
		8'd185: 32'b01110010111001001010010000000011;
		8'd186: 32'b11100011001111101101001110100001;
		8'd187: 32'b10101000110111011110000110011011;
		8'd188: 32'b01100100100100100101000100111010;
		8'd189: 32'b10010101101011100100000110111001;
		8'd190: 32'b10010111110101101010111101010011;
		8'd191: 32'b10011101000111001110001001001101;
		8'd192: 32'b11001000001001110100000110000101;
		8'd193: 32'b01010111101101111101111011001011;
		8'd194: 32'b00110101101001110000011010010100;
		8'd195: 32'b10111010001001101010111111101011;
		8'd196: 32'b10101010111011011001011010110011;
		8'd197: 32'b11100100111110111111011100110110;
		8'd198: 32'b11100001000110111011100011110011;
		8'd199: 32'b00100001001011100100001101010010;
		8'd200: 32'b01000100010010011100110111011001;
		8'd201: 32'b10010010110010001100011110101001;
		8'd202: 32'b10010101000101010000001000001001;
		8'd203: 32'b10000011110100000110101001000110;
		8'd204: 32'b01100011000101111100010111111110;
		8'd205: 32'b01010111011010110010111000000001;
		8'd206: 32'b11100111010100101111111111100011;
		8'd207: 32'b10100000011001010011101010110011;
		8'd208: 32'b11100011011100110110010011111010;
		8'd209: 32'b01111111001011011100011001010100;
		8'd210: 32'b01001001110001000110110100000100;
		8'd211: 32'b10100110001010111111001110100011;
		8'd212: 32'b11011110111110101010011101110111;
		8'd213: 32'b00110010111110010111001010101101;
		8'd214: 32'b10100001110101111000111101110101;
		8'd215: 32'b10111110000001100010100001101000;
		8'd216: 32'b11111011110000001101110110010100;
		8'd217: 32'b10001100000000001010011010010110;
		8'd218: 32'b11101110010001101101011111010010;
		8'd219: 32'b10010101010100111001110011110001;
		8'd220: 32'b00101100101011110100011110111011;
		8'd221: 32'b11100001000011010101110011010000;
		8'd222: 32'b00010011110010110110110101000101;
		8'd223: 32'b11011100110001101110001111011001;
		8'd224: 32'b00100100001110111011110000110101;
		8'd225: 32'b10010100000010100101000011011100;
		8'd226: 32'b10001110011010110101101110110010;
		8'd227: 32'b00101010010001011000110111100111;
		8'd228: 32'b11010110101001001000000000100011;
		8'd229: 32'b01010110110001011010001111010011;
		8'd230: 32'b01101001011101101000001001011101;
		8'd231: 32'b01110100111011000101111101001111;
		8'd232: 32'b11100100110001000001111101011110;
		8'd233: 32'b11101110111000011011101100110111;
		8'd234: 32'b00100011111011010001011011001011;
		8'd235: 32'b01110000001010011110100001110111;
		8'd236: 32'b01010001000110110000000101001011;
		8'd237: 32'b11100000111110111100011000000010;
		8'd238: 32'b01000101000010000010011100101010;
		8'd239: 32'b11101110001110010011100111111001;
		8'd240: 32'b11110101101010110010011001100010;
		8'd241: 32'b01000110100001110010100001001011;
		8'd242: 32'b01000011111110111001111101110001;
		8'd243: 32'b01110010011000101010110000101011;
		8'd244: 32'b10010100111011111010000011011011;
		8'd245: 32'b01011000111110111001110011111010;
		8'd246: 32'b10011100010110100010101010110001;
		8'd247: 32'b00111001110000111101111101010001;
		8'd248: 32'b00110011011010011011110011110100;
		8'd249: 32'b01111011101010111000100100100010;
		8'd250: 32'b00011101001101000110001110001100;
		8'd251: 32'b11000110001001101000110011110011;
		8'd252: 32'b00000010001011010110100010000110;
		8'd253: 32'b10010001100001011101010001010011;
		8'd254: 32'b01001011011110100001000011001001;
		8'd255: 32'b00011000110001101001101000000111;
	endcase;
	return out;
endfunction
function Bit#(32) get_msg_bit_page1(UInt#(8) counter);
	Bit#(32) out = case(counter)
		8'd0: 32'b00110101100100110011110010110010;
		8'd1: 32'b10111000101110101001011111010110;
		8'd2: 32'b01100101000111010010000110101111;
		8'd3: 32'b00011000010100001101110011100011;
		8'd4: 32'b01101101011110100010000011100011;
		8'd5: 32'b10010101010110111111000101101100;
		8'd6: 32'b00101110010000011101010001101110;
		8'd7: 32'b01111111011111110011010001111101;
		8'd8: 32'b10101100110000111001011011111110;
		8'd9: 32'b00011011010011010110001101111000;
		8'd10: 32'b01000000001001110101010011110001;
		8'd11: 32'b11111010100110100001001011001011;
		8'd12: 32'b00000100101111001111010100000111;
		8'd13: 32'b00110000100011110000100010101110;
		8'd14: 32'b11000111111010101011001001001100;
		8'd15: 32'b00011001011000100110001110000100;
		8'd16: 32'b11001100101101100101011000100001;
		8'd17: 32'b11000011010000000000000010000001;
		8'd18: 32'b01111010011110111111110101000010;
		8'd19: 32'b01001110110010001100011011000000;
		8'd20: 32'b01100110110110010000110011011000;
		8'd21: 32'b11010101011111111000100101110010;
		8'd22: 32'b10001101111110011000000010010011;
		8'd23: 32'b11111101111110100010001111010101;
		8'd24: 32'b01011101010110001110111001000111;
		8'd25: 32'b10100100100011111101101101000101;
		8'd26: 32'b00010000011000011011000010100100;
		8'd27: 32'b11110000010110101100001110010100;
		8'd28: 32'b00000000110110001000010000010100;
		8'd29: 32'b00010000011001100011001101010111;
		8'd30: 32'b00101100111011110001001000011000;
		8'd31: 32'b01110001110011100000100100111110;
		8'd32: 32'b10110011101110110100101110100011;
		8'd33: 32'b11000000011011111000010000101010;
		8'd34: 32'b01010000110100000100100110000110;
		8'd35: 32'b10100101111001010110010011001000;
		8'd36: 32'b10111101001101111100000001010001;
		8'd37: 32'b00111100101101000101111010101010;
		8'd38: 32'b11011010100001000101111111111010;
		8'd39: 32'b10101101100001001101110000111011;
		8'd40: 32'b10001110011011010110101010101010;
		8'd41: 32'b11000111111010101000001101110010;
		8'd42: 32'b11000000110011111110001000010111;
		8'd43: 32'b11111100001100000111011011001010;
		8'd44: 32'b11100101101111011110010010001000;
		8'd45: 32'b01101011111111110011011011111100;
		8'd46: 32'b01101110110001011001100000000000;
		8'd47: 32'b11010111101010010010011011100101;
		8'd48: 32'b00000000110010100111101100011010;
		8'd49: 32'b01000110001011101011110110100100;
		8'd50: 32'b10001110111111001011001110011100;
		8'd51: 32'b01000111001000001100000000110110;
		8'd52: 32'b01111110010101000001010001010011;
		8'd53: 32'b00111011110111111111100111101010;
		8'd54: 32'b10010110100000001011110111101111;
		8'd55: 32'b00100001000100010000100110000000;
		8'd56: 32'b00100100011000111111110111000111;
		8'd57: 32'b11100110101111011001111100010010;
		8'd58: 32'b00010110010111000001001110011101;
		8'd59: 32'b11101000001101011010001100000101;
		8'd60: 32'b00100100001011100111111101000011;
		8'd61: 32'b01010000001111000110011101011110;
		8'd62: 32'b01010110000011110101011000110101;
		8'd63: 32'b01100001000001110001001101111001;
		8'd64: 32'b01010111011001000111011000010100;
		8'd65: 32'b01011001100010110001111111010111;
		8'd66: 32'b11010100100010000101000111110010;
		8'd67: 32'b11010001011110100011000010010011;
		8'd68: 32'b10000010111110101111100000000100;
		8'd69: 32'b10001010111001011010011101011100;
		8'd70: 32'b01101111010010100110000110110100;
		8'd71: 32'b00100010011011001000001111001010;
		8'd72: 32'b01001010001000111000101111111001;
		8'd73: 32'b00110110010100111011000010010101;
		8'd74: 32'b11011101110111111001100101011110;
		8'd75: 32'b01010100110111110011111000100110;
		8'd76: 32'b10100101111010010101101010001001;
		8'd77: 32'b01101000111011000111110010111000;
		8'd78: 32'b00101010111110110010110110011111;
		8'd79: 32'b00111001001101110001011001110000;
		8'd80: 32'b00101101100011001110001111010011;
		8'd81: 32'b10100100010010110010000110000111;
		8'd82: 32'b01110001011000101000111011011011;
		8'd83: 32'b10100010101110000101101110011101;
		8'd84: 32'b10000011101001101111111101011111;
		8'd85: 32'b11000001111100000011000001011110;
		8'd86: 32'b01100011000011100011000110110111;
		8'd87: 32'b10011010111001001111000111110111;
		8'd88: 32'b11101100010110000101110010100111;
		8'd89: 32'b11001011001011100101110011010011;
		8'd90: 32'b00001000110000110011011111011000;
		8'd91: 32'b01001110000010000000111000001111;
		8'd92: 32'b11111001101111101101011011000010;
		8'd93: 32'b10101011101101111100001010100101;
		8'd94: 32'b00011010101010110111100000100001;
		8'd95: 32'b01000001001001000111100010111100;
		8'd96: 32'b11111010011011000111011100100011;
		8'd97: 32'b10110011111110110000011001000100;
		8'd98: 32'b10011100100010111001110101010010;
		8'd99: 32'b11000010000000111000101011001001;
		8'd100: 32'b00110111110011101100110110101010;
		8'd101: 32'b11010100101111001001110011110100;
		8'd102: 32'b01010001000000100100010101000101;
		8'd103: 32'b00110000000010101100100110010001;
		8'd104: 32'b00000001001101010001000010001001;
		8'd105: 32'b01011101111100101000100010001010;
		8'd106: 32'b01011010101000111011110000101110;
		8'd107: 32'b11010001000001110100110001000101;
		8'd108: 32'b10001001111001111000110111010011;
		8'd109: 32'b10000001110011010110101110000100;
		8'd110: 32'b01111111010100011001000011000100;
		8'd111: 32'b10001000101100101101101000111100;
		8'd112: 32'b01101001010010010110110100000001;
		8'd113: 32'b10001111011100011110001101111000;
		8'd114: 32'b11110110001111110110010101100101;
		8'd115: 32'b10011001010111000111111100001100;
		8'd116: 32'b01001111000101010000000101111111;
		8'd117: 32'b01111011011010110010111010011100;
		8'd118: 32'b01000110001001000011100000111110;
		8'd119: 32'b10101010100111111101000011000100;
		8'd120: 32'b11101100111010000011010001100100;
		8'd121: 32'b01010011110010100110001100000100;
		8'd122: 32'b11101100000000101100001110001010;
		8'd123: 32'b01101001001110011100110010101000;
		8'd124: 32'b11110101101110000101101110111101;
		8'd125: 32'b00101010011110010000100011110011;
		8'd126: 32'b10110001000000111011000101110110;
		8'd127: 32'b10111011101111100011100000110000;
		8'd128: 32'b10011010001101110001111001100101;
		8'd129: 32'b00001001011100010011101010110110;
		8'd130: 32'b01101110000111110010101011110100;
		8'd131: 32'b10010000011110001101110011110000;
		8'd132: 32'b11111001011010010011100001110000;
		8'd133: 32'b01111100101101111111010001111111;
		8'd134: 32'b00010101010101010011000010110101;
		8'd135: 32'b01100110100100000100101001001101;
		8'd136: 32'b10100100100100010010111000100010;
		8'd137: 32'b01010011100110100101010101011110;
		8'd138: 32'b01101001000100100110010111110101;
		8'd139: 32'b01001100001001111111100110011110;
		8'd140: 32'b01101010010011110010010100100100;
		8'd141: 32'b01111100001001000010101111110101;
		8'd142: 32'b00110000011011101011011100001110;
		8'd143: 32'b00011100110011101010101000100111;
		8'd144: 32'b10010110000101101111110011111110;
		8'd145: 32'b00001000010010010001001001111001;
		8'd146: 32'b11111100111110110101100010100111;
		8'd147: 32'b10101101110111001001000111011100;
		8'd148: 32'b11000101001000000111010100101110;
		8'd149: 32'b11111100111101010000010010110000;
		8'd150: 32'b11010101001100011010010001001101;
		8'd151: 32'b10010001110001001000011011001111;
		8'd152: 32'b00001011100001000110111000010011;
		8'd153: 32'b00001010011111001001110011011111;
		8'd154: 32'b10100100101010101110101001110101;
		8'd155: 32'b00110010110000111001001100100001;
		8'd156: 32'b10000000010111100110111101100110;
		8'd157: 32'b11100011111110011100011000001101;
		8'd158: 32'b00011110000001010111000010110011;
		8'd159: 32'b01101001101001011110110010000101;
		8'd160: 32'b11011111100111010001000100111011;
		8'd161: 32'b01111000111000000111000000110110;
		8'd162: 32'b01101010101101110110100010110000;
		8'd163: 32'b01011000000110111000100110010100;
		8'd164: 32'b11110000101010011101001011111100;
		8'd165: 32'b10100000001100000011001010111001;
		8'd166: 32'b01101010001011010101010110001001;
		8'd167: 32'b01101110101110001000100010111001;
		8'd168: 32'b10011110001100011000111100010100;
		8'd169: 32'b00000101100101111100001111000101;
		8'd170: 32'b10010010000010111100110101110101;
		8'd171: 32'b10001100110001110111011100001000;
		8'd172: 32'b11011010011000100110111110001101;
		8'd173: 32'b11010011110100100111100011000110;
		8'd174: 32'b00010111000010001011110010101101;
		8'd175: 32'b01111100011100010111110100010100;
		8'd176: 32'b11001101000001010111000011110001;
		8'd177: 32'b01011001001010001100100100100010;
		8'd178: 32'b00100011001001110001011011100010;
		8'd179: 32'b10111101010011111010100011001011;
		8'd180: 32'b00001111111000111010100100001111;
		8'd181: 32'b01001000011010011001001111010101;
		8'd182: 32'b11111100101101111011000111111101;
		8'd183: 32'b00011101100110010000101100000110;
		8'd184: 32'b01010010101111111110100011000100;
		8'd185: 32'b01011101011010000000010011101101;
		8'd186: 32'b11001000111111001010100000110101;
		8'd187: 32'b10101101000000100100111011001000;
		8'd188: 32'b11010011100011011101001011011011;
		8'd189: 32'b11101001101001111001100000111000;
		8'd190: 32'b01010110110100111001011100110001;
		8'd191: 32'b00101011010111000100010101101011;
		8'd192: 32'b11100011011101101111101000100011;
		8'd193: 32'b01001001000010110110110011001100;
		8'd194: 32'b01100001001010011010001010100001;
		8'd195: 32'b10101111000111111000010010010111;
		8'd196: 32'b10011000011111000001100000010000;
		8'd197: 32'b00111001011010000101011010100111;
		8'd198: 32'b01011010000001100100100110110010;
		8'd199: 32'b10011010100111000001000010110010;
		8'd200: 32'b01110011011111011100101110110110;
		8'd201: 32'b11000111011110111100110100110100;
		8'd202: 32'b00000011101110011100101101111010;
		8'd203: 32'b00111010001000110110101000100001;
		8'd204: 32'b11000110101011001001101110000010;
		8'd205: 32'b00001101010101111000010110110100;
		8'd206: 32'b11010101011001010010101110110011;
		8'd207: 32'b11111101101111110011111100000010;
		8'd208: 32'b11010000011111111110010000011111;
		8'd209: 32'b00010110101110100100100000100110;
		8'd210: 32'b00011101010101111111010100101110;
		8'd211: 32'b01000110111110001101011000000011;
		8'd212: 32'b11111110010110100010000000110101;
		8'd213: 32'b00001010101100000110101110011010;
		8'd214: 32'b00101110100101011011010110000010;
		8'd215: 32'b10100000100001011000010011100101;
		8'd216: 32'b11010111011001010011101001000011;
		8'd217: 32'b01101111011011100110100011110001;
		8'd218: 32'b00101010001001110100010100110101;
		8'd219: 32'b10001110110000111110111011100001;
		8'd220: 32'b01110101011011011111011011000000;
		8'd221: 32'b11101011110000000101110011100110;
		8'd222: 32'b00111001000101000111011110110110;
		8'd223: 32'b10100010010101101010001000111100;
		8'd224: 32'b10000000100000000001110111110110;
		8'd225: 32'b00100101011111101010110100101101;
		8'd226: 32'b11111000001000011100001010000111;
		8'd227: 32'b01111111000110010111001000110011;
		8'd228: 32'b11111101010110101001001111000001;
		8'd229: 32'b01110100101011110010001001010010;
		8'd230: 32'b00000101001000010011001110010010;
		8'd231: 32'b10000110001101100011100111111110;
		8'd232: 32'b00101010100001001110100100111011;
		8'd233: 32'b01001100010010010101100111000011;
		8'd234: 32'b11000101000010011010011011110110;
		8'd235: 32'b11000111111000000101110110111110;
		8'd236: 32'b01011101000101110100001001001101;
		8'd237: 32'b11010000111011011111011101001100;
		8'd238: 32'b01011001001001110010000011010100;
		8'd239: 32'b11010101001101110001011000110011;
		8'd240: 32'b00101010001101110111001101111010;
		8'd241: 32'b10110000101011011001101100000010;
		8'd242: 32'b10110000001010001000011010100000;
		8'd243: 32'b00101111011011010100010100100100;
		8'd244: 32'b00101011001000010110101011111011;
		8'd245: 32'b00001110111111111011100110101011;
		8'd246: 32'b11000000000110111000111100010110;
		8'd247: 32'b10000110011101101011011100101010;
		8'd248: 32'b00011100110111100110110101100001;
		8'd249: 32'b11000011001110110001100011001100;
		8'd250: 32'b00011101001100100011100011000101;
		8'd251: 32'b01000011111011100000010001010101;
		8'd252: 32'b10100011001100001100010111110101;
		8'd253: 32'b00011010000100100010011101000001;
		8'd254: 32'b01110000100011100011100100100110;
		8'd255: 32'b11010010011011010000000001100110;
	endcase;
	return out;
endfunction
function Bit#(32) get_msg_bit_page2(UInt#(8) counter);
	Bit#(32) out = case(counter)
		8'd0: 32'b11110101001101000111111101010100;
		8'd1: 32'b00011101111101010100000000101111;
		8'd2: 32'b00101000010101000001010110111000;
		8'd3: 32'b00111100000110010001111111100000;
		8'd4: 32'b11010110100011111101000110000001;
		8'd5: 32'b11001001110000110011001111001110;
		8'd6: 32'b11001001000111100001000110011101;
		8'd7: 32'b00100010101010100110101110100110;
		8'd8: 32'b01001110010000111000010010101001;
		8'd9: 32'b00110111101011010010100110010101;
		8'd10: 32'b10011101100010010001110011100000;
		8'd11: 32'b10110100101110110001001001010110;
		8'd12: 32'b01111001110100111100100101111111;
		8'd13: 32'b01101110000000100101111011100110;
		8'd14: 32'b01000111010011011011100010111001;
		8'd15: 32'b01111010110000011101000111110001;
		8'd16: 32'b00000110101000101100100011100001;
		8'd17: 32'b00010101100111011111011100000111;
		8'd18: 32'b11001110011011001110111001000110;
		8'd19: 32'b11101000100110101100110111010001;
		8'd20: 32'b10001110010111111100011000100100;
		8'd21: 32'b00001110100100100111010000110111;
		8'd22: 32'b01010101100110100011100000000101;
		8'd23: 32'b11010101010111011011110110001011;
		8'd24: 32'b01001101110100100110000111110001;
		8'd25: 32'b10010111010001001101000011100000;
		8'd26: 32'b01001101000110100110010011110001;
		8'd27: 32'b11111101000011010100000110111001;
		8'd28: 32'b10110001100101001100110001001010;
		8'd29: 32'b00101100000000101010111010000011;
		8'd30: 32'b01110100110011001110000101110111;
		8'd31: 32'b01001110010010001100101101110010;
		8'd32: 32'b11101111010000011011011101101011;
		8'd33: 32'b00110001110111010010110111101111;
		8'd34: 32'b11100111010100001001011110011110;
		8'd35: 32'b00111110010001110001111110101111;
		8'd36: 32'b11110110000001000110101000001000;
		8'd37: 32'b00101111001111010110111111100011;
		8'd38: 32'b10011101011111101010101110000110;
		8'd39: 32'b00011110010110100111111000101000;
		8'd40: 32'b00000110011111101101001101101111;
		8'd41: 32'b00001111000100111011100110101000;
		8'd42: 32'b11110100110100010101010100110100;
		8'd43: 32'b10001110101010111011000010000100;
		8'd44: 32'b01011111001001011101010001011101;
		8'd45: 32'b00001001001001101001000101001100;
		8'd46: 32'b00110010000000011111101110011101;
		8'd47: 32'b10000110010001110101110011111111;
		8'd48: 32'b01111000011110011001000011110101;
		8'd49: 32'b11011100101011111000011000000101;
		8'd50: 32'b10001100001110101111011111111010;
		8'd51: 32'b10111110011010101100000101101111;
		8'd52: 32'b00110000001100000101001001100110;
		8'd53: 32'b00101101101101100110000000100010;
		8'd54: 32'b10001011100001111000110111001101;
		8'd55: 32'b10000111111011010100000011111010;
		8'd56: 32'b01010100101010011011001010000101;
		8'd57: 32'b01100110000001011000110010101110;
		8'd58: 32'b11110010101101111000000010001011;
		8'd59: 32'b01010111010101111100110011011010;
		8'd60: 32'b10001001010111011000000100100011;
		8'd61: 32'b11110010100100001001001000100110;
		8'd62: 32'b10110000001100101101000100000010;
		8'd63: 32'b10100100101000111000010111101111;
		8'd64: 32'b10000010001101010001010101010100;
		8'd65: 32'b00000011110011101011111001011011;
		8'd66: 32'b11111010110110110100000000101110;
		8'd67: 32'b11111110011010010110101111001001;
		8'd68: 32'b00101100010111101001011001001001;
		8'd69: 32'b11110100011101011111001101010101;
		8'd70: 32'b11111100111001111001000000101000;
		8'd71: 32'b11111001100100010010101100101100;
		8'd72: 32'b11010001111110110010001010010111;
		8'd73: 32'b10001100110111001010010100110110;
		8'd74: 32'b01010000111001111010001001011011;
		8'd75: 32'b10101100110010011101011011100001;
		8'd76: 32'b01101100101100111000011001011011;
		8'd77: 32'b01011001101010110100101101011010;
		8'd78: 32'b01011100011000111000010101000000;
		8'd79: 32'b11100001111111111000110011011100;
		8'd80: 32'b10011111001101110101101010010011;
		8'd81: 32'b10110000111000101010101001011011;
		8'd82: 32'b11011110100010010111000111110100;
		8'd83: 32'b00011011101011101011101101101001;
		8'd84: 32'b01110100111001001101001111010001;
		8'd85: 32'b11001101010010101100000010000110;
		8'd86: 32'b01110111100001010111110110000100;
		8'd87: 32'b00111000001110110100001101110010;
		8'd88: 32'b10111111101110010001100001000110;
		8'd89: 32'b00000111110001100000011000111011;
		8'd90: 32'b00111111011110001010111000001010;
		8'd91: 32'b00011100100110011011011000100011;
		8'd92: 32'b00010101011010000111100101011001;
		8'd93: 32'b10100111000101010100100100011111;
		8'd94: 32'b10110101011011001011111100101110;
		8'd95: 32'b00101001010100111000101110010100;
		8'd96: 32'b11101111111111001001011110101000;
		8'd97: 32'b01001001000001000000011101011100;
		8'd98: 32'b11100011011001100111101111000010;
		8'd99: 32'b10010001101001110011111011000111;
		8'd100: 32'b00110110111111011111000101111110;
		8'd101: 32'b01001001001110011101010101110011;
		8'd102: 32'b11100001001000101001000000001001;
		8'd103: 32'b11100001101110001101110100010001;
		8'd104: 32'b01101001011000100000101111101110;
		8'd105: 32'b11110000101110111110011010010110;
		8'd106: 32'b10001110011010010111101001101101;
		8'd107: 32'b10101100001001001011101001011001;
		8'd108: 32'b10101110010001101011000111000000;
		8'd109: 32'b10011000100001110101100001001001;
		8'd110: 32'b10010101000011111110010100001101;
		8'd111: 32'b01000100010110011011110000101001;
		8'd112: 32'b00010001001000111100010110011001;
		8'd113: 32'b11010000000000100101111111100100;
		8'd114: 32'b11000011011111100001000111110000;
		8'd115: 32'b10010010101101010101000001001010;
		8'd116: 32'b01011111011101101000111111101000;
		8'd117: 32'b11000001110011101101100000100111;
		8'd118: 32'b00111001110010001000010011101010;
		8'd119: 32'b01100110111110001110100110100001;
		8'd120: 32'b01010001101011111010011100000010;
		8'd121: 32'b10100100111101100001100000111011;
		8'd122: 32'b11010001111101101110101000100111;
		8'd123: 32'b11010010010101000000011100110111;
		8'd124: 32'b01100011100000100101000010101010;
		8'd125: 32'b10000110010110111111000000110010;
		8'd126: 32'b00010001010111111001100001101111;
		8'd127: 32'b00000000101000000100111101100000;
		8'd128: 32'b10010111001011000001110101111011;
		8'd129: 32'b10001100101011111110100100111011;
		8'd130: 32'b10110100110011010000101101001011;
		8'd131: 32'b01011100011110110101111111000011;
		8'd132: 32'b00110111100100011001001001000110;
		8'd133: 32'b11111111001101010101011110010101;
		8'd134: 32'b01000100100110000110101010100000;
		8'd135: 32'b10101000110100001000111001011111;
		8'd136: 32'b01101000010101010010000001110100;
		8'd137: 32'b11100000010000010001110111100100;
		8'd138: 32'b01000101001100111100111001010001;
		8'd139: 32'b11011101100001101100110100011110;
		8'd140: 32'b10010001110110101000001011111100;
		8'd141: 32'b11011011101101101011010011111110;
		8'd142: 32'b01100001111010001111000100111001;
		8'd143: 32'b01000110011100101101011011100111;
		8'd144: 32'b11001101011100101111110100001100;
		8'd145: 32'b01100101101000000110110100000100;
		8'd146: 32'b10011000011110010101100100110111;
		8'd147: 32'b01100001001000100010010011101011;
		8'd148: 32'b11110001111111010110001000000011;
		8'd149: 32'b11011100011111100001010001000000;
		8'd150: 32'b11010101101010111100111011000101;
		8'd151: 32'b00011011101011100000001101111100;
		8'd152: 32'b00001000111010100100000001000011;
		8'd153: 32'b01100110100110010111111010111011;
		8'd154: 32'b01000000101011110010000011010100;
		8'd155: 32'b10010100011010101111011010101101;
		8'd156: 32'b00111101100000011101011011110001;
		8'd157: 32'b00100100101101000001010001110101;
		8'd158: 32'b10110011111110001100000101001110;
		8'd159: 32'b10000100111010100110011001011110;
		8'd160: 32'b11000111010000011000111101010000;
		8'd161: 32'b11011100010011001101101000101111;
		8'd162: 32'b01011101101111000101000101000001;
		8'd163: 32'b10010110000010100001000011100000;
		8'd164: 32'b10100001111001111011111110111001;
		8'd165: 32'b01101101100011001010000010110011;
		8'd166: 32'b01001101010011000010000000000010;
		8'd167: 32'b00000100010110001000001110000011;
		8'd168: 32'b10011001110000111000101010111110;
		8'd169: 32'b00011100100101110111100011100001;
		8'd170: 32'b10010011110010101001011011001011;
		8'd171: 32'b01111011000100100001011101100010;
		8'd172: 32'b10011110110111001111011000110101;
		8'd173: 32'b00010011000111011010101111010101;
		8'd174: 32'b10101011101110100010110111000110;
		8'd175: 32'b11010011100010011010001111001011;
		8'd176: 32'b10010111110100111111011011111010;
		8'd177: 32'b11110010011111011011100110100001;
		8'd178: 32'b01110101000000001110111111100000;
		8'd179: 32'b01110101100111011101110111110101;
		8'd180: 32'b01010011100011101010100101100110;
		8'd181: 32'b11010001001000011111110011100011;
		8'd182: 32'b10101000110110100001000101111001;
		8'd183: 32'b11100010001100110000000011111010;
		8'd184: 32'b10101000010110011010101011010100;
		8'd185: 32'b01000101100100011100011000011100;
		8'd186: 32'b01111011000011010100101010110111;
		8'd187: 32'b10010110000010010100101010011010;
		8'd188: 32'b00001111111011101001111010011011;
		8'd189: 32'b01010001011001100111111011111001;
		8'd190: 32'b00101011101101110100000101011100;
		8'd191: 32'b00011010111101111001010011010010;
		8'd192: 32'b11111110011110000010110011111101;
		8'd193: 32'b00101110101110100101110001010010;
		8'd194: 32'b01011100101111110101010101110011;
		8'd195: 32'b01010010001110011101101111110110;
		8'd196: 32'b10100010001000001010100100111001;
		8'd197: 32'b10100110011111110011011000001011;
		8'd198: 32'b00100010101111000011100011101001;
		8'd199: 32'b11011010111111111000001100001100;
		8'd200: 32'b10110111001001001001001010110110;
		8'd201: 32'b01101101101001111010010111110011;
		8'd202: 32'b10110110110110111111101111100110;
		8'd203: 32'b11110010110001001111101101111110;
		8'd204: 32'b11101011011101110101101001000010;
		8'd205: 32'b11000010011100101111001110001001;
		8'd206: 32'b00010011000100000100111110011111;
		8'd207: 32'b10011101011010010001001001000000;
		8'd208: 32'b10000000111101110000101000001010;
		8'd209: 32'b10011101100010001111011001011101;
		8'd210: 32'b01000110011001000011011110110011;
		8'd211: 32'b01000110001000101011001001010000;
		8'd212: 32'b10110100100100001001000101101010;
		8'd213: 32'b11001000010111100010010000111111;
		8'd214: 32'b01010001100000000111010100010110;
		8'd215: 32'b00100100101101101001100011011101;
		8'd216: 32'b11001011111101011100000011010001;
		8'd217: 32'b11111000110101101100111111101011;
		8'd218: 32'b11001011100010110011101111111101;
		8'd219: 32'b01000000100111101110010110001101;
		8'd220: 32'b11000101110010110011111010000011;
		8'd221: 32'b00000010001001010110001010011010;
		8'd222: 32'b10001110011010111101001001011110;
		8'd223: 32'b00100111100010001110101110000101;
		8'd224: 32'b10010010100111100000010110100011;
		8'd225: 32'b10110111010010101110101011000111;
		8'd226: 32'b10001110100010010000110000110110;
		8'd227: 32'b00001100011001101101011010101111;
		8'd228: 32'b10011011001011001011011110011000;
		8'd229: 32'b01001011110101110011110011001010;
		8'd230: 32'b00000010110111100100100010010111;
		8'd231: 32'b11000100101111111011000011011001;
		8'd232: 32'b11110100000001001101100001111011;
		8'd233: 32'b10100011001011011100101000111100;
		8'd234: 32'b00111011001000010010011100111010;
		8'd235: 32'b01011101111001010010000010001111;
		8'd236: 32'b01000010110010110000101011001111;
		8'd237: 32'b01001010100101100100000111101111;
		8'd238: 32'b11001101011011100000000101001101;
		8'd239: 32'b00100010011010000101111001000011;
		8'd240: 32'b00100000011101010110100010110011;
		8'd241: 32'b01001000010011101011010011110000;
		8'd242: 32'b01001000010010100001110100100010;
		8'd243: 32'b10110010101011010111000010011011;
		8'd244: 32'b01011000000101011101000110111000;
		8'd245: 32'b10110001101011101100011110000111;
		8'd246: 32'b00111110010010111001000100001000;
		8'd247: 32'b00011110000010100000111100101001;
		8'd248: 32'b10011110101110000000010010000111;
		8'd249: 32'b11000101101000001101011100101011;
		8'd250: 32'b10011011100100100000111011011011;
		8'd251: 32'b00100111001100010101100000000010;
		8'd252: 32'b01100000000101101010100100001111;
		8'd253: 32'b10110110001010000101110010101111;
		8'd254: 32'b11010001110011001111110011111100;
		8'd255: 32'b10101000100111011100111001001010;
	endcase;
	return out;
endfunction
function Bit#(32) get_msg_bit_page3(UInt#(8) counter);
	Bit#(32) out = case(counter)
		8'd0: 32'b01001110111100101100010011110011;
		8'd1: 32'b01111000111001100000100101001001;
		8'd2: 32'b00011001010100011111010110101010;
		8'd3: 32'b11001011100011001101101001011110;
		8'd4: 32'b01000101010000001011111010001110;
		8'd5: 32'b11011110110000001010000001111001;
		8'd6: 32'b01110111100010111001010001100111;
		8'd7: 32'b00001000011101011111001001010001;
		8'd8: 32'b10010110110011010110010101011000;
		8'd9: 32'b11011010011010001011001001110011;
		8'd10: 32'b00110101100101111110001100111100;
		8'd11: 32'b01000100111000001101010100010011;
		8'd12: 32'b00010101101010100111101010111011;
		8'd13: 32'b01011000101011110101111001101001;
		8'd14: 32'b10001110010101010011010010100010;
		8'd15: 32'b00111101101001001001010110001011;
		8'd16: 32'b00101000111011000101001011010000;
		8'd17: 32'b00100000000111111001110111101001;
		8'd18: 32'b01101110110110110010010001011010;
		8'd19: 32'b00010000011010011111110100001000;
		8'd20: 32'b11010010101000011111010011110011;
		8'd21: 32'b00101000100100001101110110000000;
		8'd22: 32'b01011111010100011010110111100110;
		8'd23: 32'b11011110001010000001011001001010;
		8'd24: 32'b10101000001111100010000110100100;
		8'd25: 32'b10101011110000000100000011010111;
		8'd26: 32'b11010001011010000110000101000100;
		8'd27: 32'b00110101010000001000110010001100;
		8'd28: 32'b11100000010111011010010100111110;
		8'd29: 32'b10100011110110000001001110001010;
		8'd30: 32'b10000110110101100011011111011101;
		8'd31: 32'b00000001100101110010111101110000;
		8'd32: 32'b01101110001011110100001110001101;
		8'd33: 32'b11110000011111111111000100100111;
		8'd34: 32'b10010111001000011000011111010011;
		8'd35: 32'b00010000101101000000001000101001;
		8'd36: 32'b00101010010011110101000100010000;
		8'd37: 32'b11101100000111000011101100111000;
		8'd38: 32'b11110100110101011100001111101000;
		8'd39: 32'b10001101001000011111001110011111;
		8'd40: 32'b01100110011000111000001100111010;
		8'd41: 32'b01010111111111001011100001100001;
		8'd42: 32'b11001010111010000011111010101010;
		8'd43: 32'b01101010001110000111101000010010;
		8'd44: 32'b10000101100110101101101000100111;
		8'd45: 32'b11111101110111010010011101111000;
		8'd46: 32'b01101011000011100100110111111111;
		8'd47: 32'b11001100110010010001011001101100;
		8'd48: 32'b00010101101111100110111010111010;
		8'd49: 32'b11100100101100001011100101110100;
		8'd50: 32'b00101111001111000100000001010011;
		8'd51: 32'b11010011100111101101010000011000;
		8'd52: 32'b10011010101110011001011110110100;
		8'd53: 32'b11000100101111110100101111001110;
		8'd54: 32'b11001011001110101010100101011101;
		8'd55: 32'b11011110100000110110101101000011;
		8'd56: 32'b11110000001101111011111111001111;
		8'd57: 32'b01101100011000001000000100110101;
		8'd58: 32'b01101110111111110111101011000111;
		8'd59: 32'b10101101000110011100011111101100;
		8'd60: 32'b11010111000101111110101000011010;
		8'd61: 32'b00111010010001110010000101101101;
		8'd62: 32'b10010111001111100111011001011111;
		8'd63: 32'b00110111001110001100010010101100;
		8'd64: 32'b01100100010011010010101100001101;
		8'd65: 32'b10110100010010001011101111111010;
		8'd66: 32'b10000001001011000100100110110100;
		8'd67: 32'b01110011010110100001110101101100;
		8'd68: 32'b11011110001011100100000100101000;
		8'd69: 32'b01111100001011001001110010001001;
		8'd70: 32'b10000010000101100000000000111010;
		8'd71: 32'b11001000100010101111011111100111;
		8'd72: 32'b10011100000100011011010110111101;
		8'd73: 32'b00100011011000100101011100110100;
		8'd74: 32'b01101000101111110001110100010011;
		8'd75: 32'b10101000001111111101000000001000;
		8'd76: 32'b10001100110001110010000101011101;
		8'd77: 32'b11101110101101001100111110001100;
		8'd78: 32'b10000110011110100000000011000010;
		8'd79: 32'b11111000101110101000111000101000;
		8'd80: 32'b10100000101000011000100011101011;
		8'd81: 32'b10101110001110111110101010001101;
		8'd82: 32'b01001011100101010011101100011111;
		8'd83: 32'b10111101111101001101011111110000;
		8'd84: 32'b11111011011101110100010001000111;
		8'd85: 32'b00010110010010110100111000011001;
		8'd86: 32'b10000110011100011101100100001010;
		8'd87: 32'b10000010100010000110111101010010;
		8'd88: 32'b01001110101111010100000011111000;
		8'd89: 32'b00110100101010001010100111010101;
		8'd90: 32'b11011011110110010001110000000000;
		8'd91: 32'b00100001000101111111001011111100;
		8'd92: 32'b00010010100100011011110010101010;
		8'd93: 32'b10110010010011100000011011111010;
		8'd94: 32'b11100101000000001111101010100000;
		8'd95: 32'b01001111000100100000100000110000;
		8'd96: 32'b00001000100010101111111101101111;
		8'd97: 32'b00011001101011100010101001101001;
		8'd98: 32'b11000110001101100100011111000100;
		8'd99: 32'b10010110000010110100101011010011;
		8'd100: 32'b00001111010110101100000010110101;
		8'd101: 32'b11001100010111110011100101101100;
		8'd102: 32'b10000000001111010011100010001010;
		8'd103: 32'b00101110010011000101111101000101;
		8'd104: 32'b11001100110000111100010101100110;
		8'd105: 32'b10101001111101001100001011101101;
		8'd106: 32'b01101101101000000010001100111011;
		8'd107: 32'b11101011010011010111100000001111;
		8'd108: 32'b00000110011100001011001011110111;
		8'd109: 32'b11011110000001101011010001001100;
		8'd110: 32'b00000111011100011111001111111111;
		8'd111: 32'b11000110011001000011001110001111;
		8'd112: 32'b10011111100010101110111010011101;
		8'd113: 32'b11110001110011101100111100000000;
		8'd114: 32'b01010000100100111110111010100001;
		8'd115: 32'b10000001000100100011100000001101;
		8'd116: 32'b01001100000111100100100000100110;
		8'd117: 32'b11011100011000110001011001110101;
		8'd118: 32'b10111100010100000111101001111101;
		8'd119: 32'b01011111111000001101111110110110;
		8'd120: 32'b01111001011011101111001000000000;
		8'd121: 32'b00011010010111100101110001011111;
		8'd122: 32'b11101010100011100101100111110100;
		8'd123: 32'b11101000010001001111110011001011;
		8'd124: 32'b00111100000001110000110100000010;
		8'd125: 32'b10011001100111010001001001011101;
		8'd126: 32'b00110011001110000001000001000110;
		8'd127: 32'b10011010010100101101000010101010;
		8'd128: 32'b01101110000110011001001010111110;
		8'd129: 32'b01100011000010001001010100000110;
		8'd130: 32'b01011111110001111000100001100001;
		8'd131: 32'b11101100110001000110100010111000;
		8'd132: 32'b00000011011000001100111000110001;
		8'd133: 32'b11011001100100001100011100100010;
		8'd134: 32'b11010111010110000001100010100001;
		8'd135: 32'b01111000000001101110101000010011;
		8'd136: 32'b00001110101111100110101111110010;
		8'd137: 32'b01010101101001001111010001110101;
		8'd138: 32'b11000000100011100011101011010001;
		8'd139: 32'b11111101000000110100100100011101;
		8'd140: 32'b00101100011110100111111010000101;
		8'd141: 32'b10111000101111101000100010100111;
		8'd142: 32'b01001010111010010101110001110110;
		8'd143: 32'b01111100110001000101000110100100;
		8'd144: 32'b11010000101100001000011111111010;
		8'd145: 32'b11100011011001101100010110000110;
		8'd146: 32'b01010110101010101000110110111100;
		8'd147: 32'b10010000001011000011100101011111;
		8'd148: 32'b01100000000010000010000010000010;
		8'd149: 32'b10010100000011011000100001100010;
		8'd150: 32'b01001010111110100011100001111000;
		8'd151: 32'b01000111001000111101000101011110;
		8'd152: 32'b01101111011100000010111010100010;
		8'd153: 32'b01000110111011100100001010001011;
		8'd154: 32'b01101001100100010100101001001101;
		8'd155: 32'b00001001100101100101011001110110;
		8'd156: 32'b11000110110000000000011101000111;
		8'd157: 32'b00110011010111011001011011000111;
		8'd158: 32'b10011111110011100101100010101010;
		8'd159: 32'b00010111010000010111101011110101;
		8'd160: 32'b00111110101101100011110000110010;
		8'd161: 32'b01001101111100111110100100001111;
		8'd162: 32'b11101100100101011001101000000110;
		8'd163: 32'b11011001001110011110100100000111;
		8'd164: 32'b01100100101111111111001010111001;
		8'd165: 32'b00000100101010101100100011011000;
		8'd166: 32'b01101100100000111001011110101011;
		8'd167: 32'b00111000010011111111101010010000;
		8'd168: 32'b01110101011010011011010100110101;
		8'd169: 32'b00111111110110000110110110011110;
		8'd170: 32'b00101100000001111100001111100001;
		8'd171: 32'b10101001101000111010011010101101;
		8'd172: 32'b10010111011000000110100000000001;
		8'd173: 32'b10111000000101001011111010001000;
		8'd174: 32'b11000011111011011110110010101110;
		8'd175: 32'b10010011010001110011100010001010;
		8'd176: 32'b11101110110001111111111010011100;
		8'd177: 32'b01100111011101101011010001110001;
		8'd178: 32'b10101101101011001100100111001110;
		8'd179: 32'b01011011010000110100010011001000;
		8'd180: 32'b11101001000101100101110001100111;
		8'd181: 32'b10001010111101010000100010000111;
		8'd182: 32'b01000000000101011001010001100100;
		8'd183: 32'b10111001001011001011100010100100;
		8'd184: 32'b00101011111000110100000111110100;
		8'd185: 32'b01111110111110010000100001110011;
		8'd186: 32'b11001011100000011111111100011011;
		8'd187: 32'b10000101011100001101010100100110;
		8'd188: 32'b00101101111001110100100100100111;
		8'd189: 32'b00010000011101111001101101111111;
		8'd190: 32'b10010110101100001111101110111010;
		8'd191: 32'b00101111100000000000111010001011;
	endcase;
	return out;
endfunction
function Bit#(32) get_msg_bit_page4(UInt#(7) counter);
	Bit#(32) out = case(counter)
		7'd0: 32'b01100111001101010110111111000101;
		7'd1: 32'b11101011111001110010010101100111;
		7'd2: 32'b00110111100101011011001111011110;
		7'd3: 32'b10111101100100101100111001100001;
		7'd4: 32'b01011001010011101100110110000111;
		7'd5: 32'b01000110110110101100000100100110;
		7'd6: 32'b00010011011111010000001111111100;
		7'd7: 32'b10010010100111101101000101110011;
		7'd8: 32'b11100010110110101011111000010011;
		7'd9: 32'b01111111110000011010011110100111;
		7'd10: 32'b01011110100100000100001001010011;
		7'd11: 32'b10011100011000100010010110001110;
		7'd12: 32'b11100010010101001110011100010000;
		7'd13: 32'b01111001101001100100100011010010;
		7'd14: 32'b10010010100000111100111111010101;
		7'd15: 32'b00100000011101011110011111100000;
		7'd16: 32'b00110000100000001111001000111101;
		7'd17: 32'b00100100011100111101111111101000;
		7'd18: 32'b01010111111010010010011011111100;
		7'd19: 32'b00001000000101101001101110010111;
		7'd20: 32'b01011110111010011100010000101001;
		7'd21: 32'b00010010010110110101110001100100;
		7'd22: 32'b10010101000110000010011011000001;
		7'd23: 32'b10000000111110101110101001011110;
		7'd24: 32'b00010001000111011110101000001000;
		7'd25: 32'b01000000100010101110111000110111;
		7'd26: 32'b01011000100101001001001010111100;
		7'd27: 32'b11010110111011111100000111000001;
		7'd28: 32'b10001001001010111001111001110111;
		7'd29: 32'b01010011110110110101001100010110;
		7'd30: 32'b10010011110001110111011100011011;
		7'd31: 32'b01101001001000110001001101100010;
		7'd32: 32'b00011101011010110100111000100001;
		7'd33: 32'b10000110101010101111101101011010;
		7'd34: 32'b11011111000101101011100011100001;
		7'd35: 32'b11001111011111010000000110001100;
		7'd36: 32'b00000011100100011010010111111100;
		7'd37: 32'b10010100010001011101110000011010;
		7'd38: 32'b10000101100110010101110111111101;
		7'd39: 32'b10111110001101101001000010010000;
		7'd40: 32'b01001100000011001110111101000111;
		7'd41: 32'b11111100001010111111101100110111;
		7'd42: 32'b11000110110111011000000101000110;
		7'd43: 32'b00010001100010100011001000111000;
		7'd44: 32'b11000100010111001000010010011111;
		7'd45: 32'b01101110010111111101011000111000;
		7'd46: 32'b01001100001101111011100000000111;
		7'd47: 32'b11110101111110010011111011000011;
		7'd48: 32'b01001011101011011111110001001001;
		7'd49: 32'b10110001010100110110011011010111;
		7'd50: 32'b00010100111001000111111011001110;
		7'd51: 32'b10101101011000101101100011110111;
		7'd52: 32'b01011100101011100111101001101110;
		7'd53: 32'b00100100100000001011000011111110;
		7'd54: 32'b10110100001110000111010001001001;
		7'd55: 32'b00111111010000111000111010101001;
		7'd56: 32'b10101110010010010011101001101001;
		7'd57: 32'b11101010001001101010110100101110;
		7'd58: 32'b11010010100111010010101111011100;
		7'd59: 32'b01001010110000110000101110001110;
		7'd60: 32'b11101001011110011001100000101000;
		7'd61: 32'b10101101001111101011000111001011;
		7'd62: 32'b00011101111010111110001000010111;
		7'd63: 32'b00011110000010010100001100000011;
		7'd64: 32'b01111101010110101010010001010101;
		7'd65: 32'b01000001001010000101011111011100;
		7'd66: 32'b11000110111001111111001011101011;
		7'd67: 32'b00110011101000101011100111111100;
		7'd68: 32'b10011110100101010011110110011110;
		7'd69: 32'b11000001010000001000100111111010;
		7'd70: 32'b10110100111110111110100000110110;
		7'd71: 32'b01110101010101101100100000100100;
		7'd72: 32'b10000111000100001011101000010111;
		7'd73: 32'b00111011011010011001010110111001;
		7'd74: 32'b00011110110111010101101010110111;
		7'd75: 32'b11011110001110010101000100001011;
		7'd76: 32'b11010100100101001001011000010100;
		7'd77: 32'b11010110110111110100110011001111;
		7'd78: 32'b00011110010111100000000001111101;
		7'd79: 32'b11100010101010110010010100000011;
		7'd80: 32'b01011001100010010000100001110011;
		7'd81: 32'b11100010101100101111001110010011;
		7'd82: 32'b10110010010101011011010101000001;
		7'd83: 32'b00100111100100001101000000000110;
		7'd84: 32'b00110110111001001010001100010101;
		7'd85: 32'b01100010010101001100100000000111;
		7'd86: 32'b01000010101110010011001010101000;
		7'd87: 32'b11000000001101110010100111011110;
		7'd88: 32'b00010011110101111011100101010000;
		7'd89: 32'b10101010101100010110010100011110;
		7'd90: 32'b10001001000001010111101101110001;
		7'd91: 32'b10010010010000001011001010100010;
		7'd92: 32'b10001011111010111110011100101100;
		7'd93: 32'b01001101110100011100011011001001;
		7'd94: 32'b00010010101101101101111000011101;
		7'd95: 32'b10100001100011100111011110010110;
		7'd96: 32'b00100101101111001010001110000001;
		7'd97: 32'b10111000111000111111100110101001;
		7'd98: 32'b01110001100010001010111100001101;
		7'd99: 32'b11100111001000011011111100100111;
		7'd100: 32'b01011111001101100111111110100010;
		7'd101: 32'b11000111011101010100011011101101;
		7'd102: 32'b01111100110100000100010100110011;
		7'd103: 32'b00000010110010001110000000101100;
		7'd104: 32'b11101000111110100111110001111100;
		7'd105: 32'b01110101101011111111111001100011;
		7'd106: 32'b11111000001000101111010101101100;
		7'd107: 32'b11011101000111100000010001011000;
		7'd108: 32'b00001011101100101111100100111001;
		7'd109: 32'b10111001010000011001000000110110;
		7'd110: 32'b00000111000010101001101001000100;
		7'd111: 32'b01111101011001001101001010111110;
		7'd112: 32'b11000110000110101010111000011110;
		7'd113: 32'b00010100111010100101011101000011;
		7'd114: 32'b10011011101001101001100101110110;
		7'd115: 32'b11001110011000101010110000110111;
		7'd116: 32'b01011101101111000100101110110000;
		7'd117: 32'b00000111011111001110001101010010;
		7'd118: 32'b10101100101010000100111111101101;
		7'd119: 32'b01101010110100100111101001100110;
		7'd120: 32'b01010110110111101111010000001111;
		7'd121: 32'b10110111000111011001000101111010;
		7'd122: 32'b11001111001001111111001000010100;
		7'd123: 32'b10100010000011110010001001101010;
		7'd124: 32'b10001110010000101110110010001010;
		7'd125: 32'b10100010100111111110010000110011;
		7'd126: 32'b11100000010001101000100110000010;
		7'd127: 32'b01100011100111010010001100011110;
	endcase;
	return out;
endfunction
function Bit#(32) get_msg_bit_page5(UInt#(7) counter);
	Bit#(32) out = case(counter)
		7'd0: 32'b01101010100010011100001101101000;
		7'd1: 32'b11010001011110110010010010011001;
		7'd2: 32'b10000110011001000001000000001111;
		7'd3: 32'b11010110110001000101011110100011;
		7'd4: 32'b00000110010100111000100011011000;
		7'd5: 32'b00000001110101101011010011101001;
		7'd6: 32'b11100100011111110111100111111100;
		7'd7: 32'b10000111011110100001110011000010;
		7'd8: 32'b01111100010011011000101110100101;
		7'd9: 32'b10001101110110000110110110010000;
		7'd10: 32'b11111100101101111010110111000010;
		7'd11: 32'b10101011001101101100010000110110;
		7'd12: 32'b10111111111001111100000101001101;
		7'd13: 32'b10101110111110101101111111000011;
		7'd14: 32'b11110001000000111110001101101001;
		7'd15: 32'b10001110101101100000111010101010;
		7'd16: 32'b11110111101101010111011110101010;
		7'd17: 32'b11101101001101010010000100011011;
		7'd18: 32'b00111111100110001011100100000101;
		7'd19: 32'b01000101100000011011000100000101;
		7'd20: 32'b00001001110010000100010010100100;
		7'd21: 32'b11111000101111011111011111000110;
		7'd22: 32'b11110110001010101101101000111010;
		7'd23: 32'b10010100000100001001111001101000;
		7'd24: 32'b01101111101000110111001001100111;
		7'd25: 32'b11100100110001011001100011101110;
		7'd26: 32'b01011001011000110111011010011110;
		7'd27: 32'b10011101110111110000110101110111;
		7'd28: 32'b01100001110011110111000101110100;
		7'd29: 32'b11001010110000011001011110111010;
		7'd30: 32'b11111111000111101011101110011110;
		7'd31: 32'b01001010110100011011001000010100;
		7'd32: 32'b10111011000001100100111011101101;
		7'd33: 32'b01010110110010010100100111111011;
		7'd34: 32'b11010111111001100100000101111111;
		7'd35: 32'b11110111011011000100100010100110;
		7'd36: 32'b11011111001000010100001100000110;
		7'd37: 32'b11101111010110111111110111100001;
		7'd38: 32'b00110101011110101000110100010100;
		7'd39: 32'b01111101010100110001110110000001;
		7'd40: 32'b10000101001111111000000001101100;
		7'd41: 32'b00011111000000100111001101000110;
		7'd42: 32'b10101011100010001110100010111010;
		7'd43: 32'b00000110001111011110001011101001;
		7'd44: 32'b01001100111011000110110000110100;
		7'd45: 32'b01111111001101010101100101110010;
		7'd46: 32'b10110010000001010000100100110000;
		7'd47: 32'b00110100111110011101110100010011;
		7'd48: 32'b11010000110100010100110110111011;
		7'd49: 32'b00011111101000000010011110100101;
		7'd50: 32'b10001010000001010110001011011110;
		7'd51: 32'b01101110101100000000110010110111;
		7'd52: 32'b00101100111011001010001101000100;
		7'd53: 32'b00000001110111110000011101000001;
		7'd54: 32'b00101100100100010010111000001010;
		7'd55: 32'b01011100001001100101110111011000;
		7'd56: 32'b10111101001110000000011100000101;
		7'd57: 32'b01101110010011101000101011011101;
		7'd58: 32'b01011100010111010101100100101001;
		7'd59: 32'b10111011110000110111101001010100;
		7'd60: 32'b11001010001000010001101011010001;
		7'd61: 32'b10100110001101110111001001010001;
		7'd62: 32'b11110100101001011011101110001110;
		7'd63: 32'b11010100001011000011000100000001;
		7'd64: 32'b11111011110011000100000110000001;
		7'd65: 32'b10011001110011011101000111111111;
		7'd66: 32'b01000010000101001110110110010001;
		7'd67: 32'b10010110101000110100101100110101;
		7'd68: 32'b10111000100111111000100000111000;
		7'd69: 32'b11011110010000100111010100011001;
		7'd70: 32'b01000101010001011000000001110101;
		7'd71: 32'b00011101100100010101110000000110;
		7'd72: 32'b01010111111101101111100101111000;
		7'd73: 32'b11010111111101111010100110101010;
		7'd74: 32'b00101001010100000010011100011101;
		7'd75: 32'b11011111110111101001010011100101;
		7'd76: 32'b01000110110110101000101011011001;
		7'd77: 32'b00101001011001101100010111111000;
		7'd78: 32'b11010011111100110000111101111111;
		7'd79: 32'b11110011010100010000101000110110;
		7'd80: 32'b01010001010001000011001100101111;
		7'd81: 32'b01001110001100111101001001001111;
		7'd82: 32'b00100010001001011100000001010011;
		7'd83: 32'b01011010101101101011010010000100;
		7'd84: 32'b01000000101011111001010001001100;
		7'd85: 32'b00000111111010110011100000001110;
		7'd86: 32'b00101001110110011100010111001010;
		7'd87: 32'b00011010101010100011100101110111;
		7'd88: 32'b11111000011110110000110100101111;
		7'd89: 32'b01111111010100011100100011000100;
		7'd90: 32'b01001111110101101110111010100100;
		7'd91: 32'b11110110000010000110001000111100;
		7'd92: 32'b00111100011101010110100101100111;
		7'd93: 32'b01000010110011001101011101001011;
		7'd94: 32'b10111001001111000111000110111011;
		7'd95: 32'b11110001000100100011111110000111;
		7'd96: 32'b11101111101110011111110010000101;
		7'd97: 32'b00100010110100100000111000111011;
		7'd98: 32'b00010100000100010101011010010100;
		7'd99: 32'b01010001111000110110111101101001;
		7'd100: 32'b00110101100100011001101101101101;
		7'd101: 32'b00010000101010001100001100000000;
		7'd102: 32'b10001110000001010111100111001111;
		7'd103: 32'b00111100010101001000101001100001;
		7'd104: 32'b00011101101110001101000011101000;
		7'd105: 32'b01011001001000110110100011000110;
		7'd106: 32'b11101000010111011001001011000111;
		7'd107: 32'b01001111000000011010011110010100;
		7'd108: 32'b00000110001110001100011011100011;
		7'd109: 32'b00001010000101011101011000101011;
		7'd110: 32'b11100111001110010010101101110110;
		7'd111: 32'b00000100111010110000101000010111;
		7'd112: 32'b00110000000110110100110010000101;
		7'd113: 32'b00000010101000010100110101110000;
		7'd114: 32'b00001101111100101110001011010110;
		7'd115: 32'b10001010010110001000100001011110;
		7'd116: 32'b00111111100110110101111110001000;
		7'd117: 32'b11011111001001001101111100010101;
		7'd118: 32'b01110111101110010011110011001011;
		7'd119: 32'b01110000001111001101001010111011;
		7'd120: 32'b11100101001001011011100001111001;
		7'd121: 32'b10001011100000010101001110011111;
		7'd122: 32'b01110111101000001101101001100111;
		7'd123: 32'b00101010100101000111011111000000;
		7'd124: 32'b01101110011001110100001010001000;
		7'd125: 32'b10011001011001100011011110100110;
		7'd126: 32'b10111010111100101111100100101110;
		7'd127: 32'b00011110111001100001111010011100;
	endcase;
	return out;
endfunction
function Bit#(32) get_msg_bit_page6(UInt#(6) counter);
	Bit#(32) out = case(counter)
		6'd0: 32'b01111011110100010010111000001111;
		6'd1: 32'b10000011000011010010110000100011;
		6'd2: 32'b01000001001110011110111011100100;
		6'd3: 32'b01101001101111111101100111100011;
		6'd4: 32'b10110110101001101010110110010010;
		6'd5: 32'b01000010101101111101000111011010;
		6'd6: 32'b11101100101100010111010111110111;
		6'd7: 32'b00011100110100001000000100011111;
		6'd8: 32'b10111011001111100010100111101000;
		6'd9: 32'b00011100111011011001011101000111;
		6'd10: 32'b01010101010101000111000111101111;
		6'd11: 32'b11101101110111010001101001101010;
		6'd12: 32'b00110101100100111011101100100100;
		6'd13: 32'b00101101110101111001011000001010;
		6'd14: 32'b00101101100110100010000001010111;
		6'd15: 32'b00000110000100000010100100001010;
		6'd16: 32'b10011000101110001100011000100101;
		6'd17: 32'b11010010010001111100101101101010;
		6'd18: 32'b01110001000000101101000000111001;
		6'd19: 32'b00010101010010111001001001001100;
		6'd20: 32'b11000011111101011111100100101100;
		6'd21: 32'b10011100100000000010001111101011;
		6'd22: 32'b11001111100100000011000001111111;
		6'd23: 32'b11110101011001101111111000100110;
		6'd24: 32'b11000110000011111010100100010000;
		6'd25: 32'b11000111111100000101010111011111;
		6'd26: 32'b01101100111110100000010010110110;
		6'd27: 32'b00011011000101100111110010100110;
		6'd28: 32'b01011100111110010111101111011101;
		6'd29: 32'b00001001010011110111111100110101;
		6'd30: 32'b11001101001001001110011000111001;
		6'd31: 32'b01110100110011001001101110001001;
		6'd32: 32'b11111011010011011101000100100101;
		6'd33: 32'b10111001000100101101111011011001;
		6'd34: 32'b10001100010111010000000110001110;
		6'd35: 32'b00000111101111001100100000000010;
		6'd36: 32'b01001111010111100001010111000101;
		6'd37: 32'b00101110001000001101010101110101;
		6'd38: 32'b00001110100001110110110000011010;
		6'd39: 32'b00100100000011100001001010000010;
		6'd40: 32'b01011010101011000001101101100110;
		6'd41: 32'b00011001111111000100110101011000;
		6'd42: 32'b11011011101101001111010000010111;
		6'd43: 32'b01011100011001000001001110001100;
		6'd44: 32'b10010001001110100001011000111100;
		6'd45: 32'b11111110101001000100001011111100;
		6'd46: 32'b01010101000001100000100011010001;
		6'd47: 32'b10101101100000110001000101011001;
		6'd48: 32'b10010011101011101100000111001100;
		6'd49: 32'b10001111000000010010110111100000;
		6'd50: 32'b01011100011000111111111011001101;
		6'd51: 32'b10111110111010000000101011000000;
		6'd52: 32'b10100010111001011110010000000111;
		6'd53: 32'b10011110101010010101101011010010;
		6'd54: 32'b00011101100101011111010011101011;
		6'd55: 32'b01101111111010110000110111110001;
		6'd56: 32'b11000111011001111100010111110110;
		6'd57: 32'b00000001110101111100110001110010;
		6'd58: 32'b10111000001110000001010001011001;
		6'd59: 32'b11111001011001000101000011001100;
		6'd60: 32'b10100111000011100001000010011000;
		6'd61: 32'b10111111100101010111001111001101;
		6'd62: 32'b11001010101001001010000101010010;
		6'd63: 32'b00010111000111111111011010101110;
	endcase;
	return out;
endfunction
