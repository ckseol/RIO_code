function Bit#(64) get_output(UInt#(8) counter, UInt#(3) page_num);
	Bit#(64) enc_output = case (page_num)
		3'd0: get_output_page0(counter);
		3'd1: get_output_page1(counter);
		3'd2: get_output_page2(counter);
		3'd3: get_output_page3(counter);
		3'd4: get_output_page4(counter);
		3'd5: get_output_page5(counter);
		3'd6: get_output_page6(counter);
	endcase;
	return enc_output;
endfunction

function Bit#(64) get_output_page0(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b0000000000001000000111000000000000000000000100000000000001100000;
		8'd1: 64'b0000000000000000000001000000100000000100001000010010000000000100;
		8'd2: 64'b0000000100000000000000000000001000110000000000100000000100000000;
		8'd3: 64'b0001000000000000011000000001000000010000000000000000000000010010;
		8'd4: 64'b0000000000000100000000000110000001000000000000000000001000000100;
		8'd5: 64'b0000000000100000100000100100000001110000000000000101000001000000;
		8'd6: 64'b0001100000000000000000000000000001001000000000000000001100000000;
		8'd7: 64'b0000000101000001010000000000000000000000000010000000000100000000;
		8'd8: 64'b0000010000001000000100000000000000100001000101000010101100001000;
		8'd9: 64'b0000100000000000000000000000000000000000000000000000001100000000;
		8'd10: 64'b0000000001000000010000100010101000000000000000001000000011100000;
		8'd11: 64'b0000000010000000010000000000001000000100000000000010000000000100;
		8'd12: 64'b0000000000000010100010000000011100000000010000000000000000000100;
		8'd13: 64'b0001100001000000000001000000000000000000000000000000000000000001;
		8'd14: 64'b0000000000000000000010000100000000000000000100000000010000000000;
		8'd15: 64'b0000010000000000001010000000000000010000000010010000000001100000;
		8'd16: 64'b0100000000000000100000000000000000000000000000001000010001000000;
		8'd17: 64'b0000001100000000000000000000000000000001000001001000000000000001;
		8'd18: 64'b0000000000000000000000110000000001010001000100000000001000000000;
		8'd19: 64'b0000100000000001000000001001001000000000010000010000001000000100;
		8'd20: 64'b0010000000000000000100000100001000000000000010000000000000000000;
		8'd21: 64'b0000000001000000100000000100000000000000000000000010000000000000;
		8'd22: 64'b0000000000000000010000000000100010000000000100000000000000000011;
		8'd23: 64'b0000000000001000000000000011000000100000001000010000000001010100;
		8'd24: 64'b0000100000000000100000000000000100000000001000000000010010100000;
		8'd25: 64'b0000000000000000000000001011000000000010000001010001000000000000;
		8'd26: 64'b0000000001000101100000000000000000001000001000000000000000000000;
		8'd27: 64'b0100000001000100010001000000000000000000010000000010000001000000;
		8'd28: 64'b0000100000000000000000000000010001000000100000000000000000000000;
		8'd29: 64'b0001000010000010000001000000000000000000000000000000000000001000;
		8'd30: 64'b0001000100000000000000010001000000000000000000000000000000000000;
		8'd31: 64'b0000000000000100000000001001000000100000000000000000000000000011;
		8'd32: 64'b0101000100001000000000001100000000110010010001110000000000000000;
		8'd33: 64'b0001000000000001001001000000000000100100000001000000100000000000;
		8'd34: 64'b0000100000000001000001110000000000000001000000000000001000000000;
		8'd35: 64'b0000000100000011000000000000000110000001000000000000001000001000;
		8'd36: 64'b1000000000000000000000101000000000000001000000000010000000000000;
		8'd37: 64'b0000000000000000000000000100000000000000100000000010010100000000;
		8'd38: 64'b1001100000000000000000000100000000000000000000000000000000000010;
		8'd39: 64'b0000000000001000000000000000000000010001000011001100000000000000;
		8'd40: 64'b0101001000000000000000000000000100101010000000000010010010010000;
		8'd41: 64'b0000100100000000000000000001000000001010000000000000000000000000;
		8'd42: 64'b0000000000000100000000000000001010000000000000000100010000000000;
		8'd43: 64'b1001010000000000101000000000000000001001001000000000000000000000;
		8'd44: 64'b0100000000000000000000100000001100000000000010000000000010000010;
		8'd45: 64'b0100000000000110000001010000000001000000010000100001000000000010;
		8'd46: 64'b0000000000000000000000000000001000000100001000001000001001000000;
		8'd47: 64'b0000000001000000000000000000000100000100000000000000000000000000;
		8'd48: 64'b0000001001001000101000000000000000000000000100010010000000001000;
		8'd49: 64'b0010000000000000000000100010000100000000000000010000000000000000;
		8'd50: 64'b0001000000011000010100000010000000100000000011000000000000000000;
		8'd51: 64'b0000010000000000001000000000000001000000000000010000100110000000;
		8'd52: 64'b0000010000000000100000100000000100000000001000010100000001000001;
		8'd53: 64'b0000100010000001000000000000000001000000000000000000100100100100;
		8'd54: 64'b0000000010000000000000000110001000000100000000100000000000000000;
		8'd55: 64'b0000010011000000000000000000000000000000000100000000000000100101;
		8'd56: 64'b1100000001000000001010000000000000000000000001000000000000000000;
		8'd57: 64'b0000000010001000000000000000000000001010000000000010000100000000;
		8'd58: 64'b0000000011000000000000000100000000000100000000000000000000100100;
		8'd59: 64'b0010001000000000000000000000000000000000000001000010000100010010;
		8'd60: 64'b1010000000000111011100000000010000010000000010000000000000001000;
		8'd61: 64'b0000100000000000000000000011000000100100001000000000010000010100;
		8'd62: 64'b0000001000000000000000000100000000000000001000000001000000010000;
		8'd63: 64'b0000000000000000000100000000110100000000000000000000000001000000;
		8'd64: 64'b0000010000000000001000000001001000100000100000000000000000000000;
		8'd65: 64'b0000000000000000001000000000000000000000000000000100000000000000;
		8'd66: 64'b0100000011000010000110000001000000000000000000010000000010000100;
		8'd67: 64'b0000100000100000000010100000000000000010000000000000000000000000;
		8'd68: 64'b0000000000000100000001001000000000000000010010011000000000000000;
		8'd69: 64'b0001000000000001000000000000000000000000000000001001000000000000;
		8'd70: 64'b0000010010010000000000000000000000000000010100010000000000100000;
		8'd71: 64'b0010000000000110000000000000100000000000000001000000000000000100;
		8'd72: 64'b0000001000000010100000001000000000001000001000000000000000000000;
		8'd73: 64'b0000000000000000000000000100010101000000010000100000001000000011;
		8'd74: 64'b0000001011000000000010000000001010000010000100000000000010000100;
		8'd75: 64'b0000000000001000000000000000100000000000000100000000000001001000;
		8'd76: 64'b0000100010010000000000000001000000000000000001000000010000100010;
		8'd77: 64'b0001000000000001000000000000001000101100000100000000000000000000;
		8'd78: 64'b0000000000000000010000000100000000000000100010001100010000000100;
		8'd79: 64'b1000010010000000100010000000000000000000000010110000000000000000;
		8'd80: 64'b0000000000010000000001000001010000000100000100000010000000000000;
		8'd81: 64'b1000000000100000010000000000000001000000010000000010000000000001;
		8'd82: 64'b0100000000100000000000001001001000010000100000000000000000000000;
		8'd83: 64'b0000000010000011100010000000000000000000000000000000000100100000;
		8'd84: 64'b0100000000000000100010010000000100000000010000000000000010001100;
		8'd85: 64'b0000000000000000000000000010000000000000110001000000011000100000;
		8'd86: 64'b0000010000000000001000000000000000001001000000010011010100001000;
		8'd87: 64'b1001000000000000100000011000000000000000010011000000000000000000;
		8'd88: 64'b0000000000001010000010010000010000000000100000000000100000000000;
		8'd89: 64'b0000000000010000000000000101000000001000110000001000000000000000;
		8'd90: 64'b1000010010110100000000000000000000000001000000000010001101010100;
		8'd91: 64'b0000010000000001010000000000000000000010100000000000000000000000;
		8'd92: 64'b0000000110000000001000000000000000110000000000000000000000000001;
		8'd93: 64'b0010100000000000000000000010000000001100001000000000001001000000;
		8'd94: 64'b0001000000011010000000010000000000010001000100000000100000000010;
		8'd95: 64'b0001000100000001000000000010010000010000001000000000000000000010;
		8'd96: 64'b0010000100000010000000000000000000010000010100000001000010010000;
		8'd97: 64'b0000110000000000000000000000001001000100001000000000000000000001;
		8'd98: 64'b0000000000101000000000010110000000000000000000000100010000000000;
		8'd99: 64'b1000000000000000100000000100011000000100100001000100000100000010;
		8'd100: 64'b0000000000001000100000000000100000010000000000000101010000000000;
		8'd101: 64'b0010000010000100000011000100000000000000001001010000000000000000;
		8'd102: 64'b0000001000010000000100100000010001000000000110000001000010000000;
		8'd103: 64'b0100000000000000000100100000000000000000000000000100000100010000;
		8'd104: 64'b0000011000000010000101000000000000100000000000100000000100000000;
		8'd105: 64'b0000000000000000010010111110000000000110100000000101000000000000;
		8'd106: 64'b0100001100010001000000000100000000010000000000000100000100000000;
		8'd107: 64'b0100000100000001000010000000100000010000000001000000000000000000;
		8'd108: 64'b0000100001000000000001000000000001000000001000100000000000001000;
		8'd109: 64'b0010000000000000000010000000010000000000001000000100000000000010;
		8'd110: 64'b0000000000000011000000000000110000001000101100000000000000000000;
		8'd111: 64'b0001101010000000000000010000000000000000000000100011000100100010;
		8'd112: 64'b0000000000000100100000000000010000000000000100000010110000000011;
		8'd113: 64'b1001000000000001000100000000000000000000000001000000000000010010;
		8'd114: 64'b1001100000000000000000000000100100101000000000000000000000010001;
		8'd115: 64'b0000000110000000000000000000000000100001000000000001000000000000;
		8'd116: 64'b0000000000100001000000010000000000000001000100000000110000000000;
		8'd117: 64'b0000000100100100001010000000000001000000010001000000000100000100;
		8'd118: 64'b0110000000000001000000000000100000010000100000000000000000000000;
		8'd119: 64'b0100000000010010000000010000001010000100000010100000001010000000;
		8'd120: 64'b0000000000010011000000000000010000100010001000000100010000000001;
		8'd121: 64'b0011001011000100010000000000000000000000000000000000000000000000;
		8'd122: 64'b0000000000000000000000000000100000000000000000000000000000000100;
		8'd123: 64'b0100000000100000000100000000000000000000000010000010000000100010;
		8'd124: 64'b0000100000000010000000001010000000000000000000000000000000000000;
		8'd125: 64'b0000000000001000000000000000000000101000010001000000010000100000;
		8'd126: 64'b0000000000011010000000000000001001000000000010000000000000000001;
		8'd127: 64'b0000010000000000001010000000000100000000000000000000000000000001;
		8'd128: 64'b0000000000000000000010000000000100010000000001001000100000010010;
		8'd129: 64'b1000000000010010100000000101000000001000001000000000000000000000;
		8'd130: 64'b0000000100001000000000000001100100000000000000000001011000010100;
		8'd131: 64'b0101000001000000001110000000000010000000000000000000101000000000;
		8'd132: 64'b0010000000101000000000001010000000010001100000001110000100000000;
		8'd133: 64'b0000101000100000001010100000100000000001000010000000000000000000;
		8'd134: 64'b0000000010001000000000100110000000000000001000000100000001000000;
		8'd135: 64'b0000000000000000000000100010000000100000000000000010000000000000;
		8'd136: 64'b0010000010000000000000001000000001000000100000000010010000000000;
		8'd137: 64'b0000011100000000001001010010001000010000000101000000000100000000;
		8'd138: 64'b0001000100000100001100000000110000001100000000010100000001000100;
		8'd139: 64'b0000000010000001001010100100000000000000001000000100100000000000;
		8'd140: 64'b0000000000000000000000010000000100000000100000100000101000010000;
		8'd141: 64'b0000000000100000000010001000001010010000001100000010000100000001;
		8'd142: 64'b0100101000010000000000000001101010000000000000000000000000000001;
		8'd143: 64'b0100000001000000000000001000001000001000001000110000000000000001;
		8'd144: 64'b1000000000001100000000000100100000000001000000000000000000000000;
		8'd145: 64'b0010000010000100000001000101010000000010000000000100001001100000;
		8'd146: 64'b0000010001000000010000000100000000100000000101000000000000000100;
		8'd147: 64'b0000000000000000100000000000001100000011000000001100000010000000;
		8'd148: 64'b0000011000000000000100000000000000000000001000000000001000000100;
		8'd149: 64'b0000000000000000000000010101011000000000000000000000000001000010;
		8'd150: 64'b1000100010000000100000000000001100000000010100000000000010000000;
		8'd151: 64'b0100000000010001100101000000000000000000000000000010000001000000;
		8'd152: 64'b0000100000000000101010000000001010100100000000000000000000000000;
		8'd153: 64'b0100000010000000100100001000000000001000001000000000000000100000;
		8'd154: 64'b0000010000000000000010000100000000000000000001000000010000001110;
		8'd155: 64'b0000100000000010000001000000000000010000000001000000000000000000;
		8'd156: 64'b0000000100011001000000010000000000001000000000000000000000001010;
		8'd157: 64'b0010000100000000110100000111000010000000000000000000000000000000;
		8'd158: 64'b0000000000000000000000000000000001100000000010000000000000010010;
		8'd159: 64'b0000100001000000000000100000000000100000001000000000000001000000;
		8'd160: 64'b0000010000000010000000000000000000000000000001000000000000001000;
		8'd161: 64'b0000000000000000100000000010000000100100000000000000000000001000;
		8'd162: 64'b0100011011001000000101001100000000100000000000000100100100100000;
		8'd163: 64'b1110000000010000100001000010100000000000000100000000000000100000;
		8'd164: 64'b0000000000000001000100010000101000000000000000010010000110000000;
		8'd165: 64'b0000010000000100100010100001000100101100000001010000000000000000;
		8'd166: 64'b0000010000000001000000000000010000000000001001000010000100100000;
		8'd167: 64'b0010000010000000000000000000000111000000000000000000000001000000;
		8'd168: 64'b0000001000001000010001000000000000100000000000000000000001000000;
		8'd169: 64'b0100000000000000010100000000000000000000100000000100000010000001;
		8'd170: 64'b0000000000000100000000001000001100000000000010000000000101000000;
		8'd171: 64'b0000000010000000000000000010011000000000000010000000000000000000;
		8'd172: 64'b0010000000000101001000000001000000000001000000000010000001010000;
		8'd173: 64'b0001010001000000000000000000001001000000000000000000000000000000;
		8'd174: 64'b0000000100000000000000000000000000000000000011010100100000000000;
		8'd175: 64'b1010000010010000001000000000000000000000000000001000000000000010;
		8'd176: 64'b0010000000010101001010000000000100000101000000000010000000100000;
		8'd177: 64'b0010100010000000000001000001000000010000000001000000100010000100;
		8'd178: 64'b0000001010000000001000000000000000000000000000000000000000000000;
		8'd179: 64'b0000000000000000000000001000000100001000101000000010000001000010;
		8'd180: 64'b0010000000000000000000000000000000000000000010000000010000000010;
		8'd181: 64'b0001000010010000000000000100000010000001000000100010000000000000;
		8'd182: 64'b0000000010011000000010101000000000101001001100100000000000000000;
		8'd183: 64'b0010000010000000000000000000000000000000001101000000000110000100;
		8'd184: 64'b0010000100100000000001000000000001000010000000000000000010000000;
		8'd185: 64'b0000000000000001001000000000000001001000000000000001000000000100;
		8'd186: 64'b0000000001100010000000001001001000000000000100000100000101000000;
		8'd187: 64'b1000000001000000000000000000000001001100000000010001000000000010;
		8'd188: 64'b0000001000000000000011000001000000000000000000100000001000000000;
		8'd189: 64'b0000000000000011000000000000010000000000000000001000000000100110;
		8'd190: 64'b0000000000010000000000000110000001000100001101000000000000000001;
		8'd191: 64'b0100000001101000000001100000000000010010000000100001100000000000;
		8'd192: 64'b0000000000000001001000100000001000000000000000100101010000000000;
		8'd193: 64'b0101000001100100000000000000000000000110000000000001000000000001;
		8'd194: 64'b1000000000000100000100000000000000000101100001010001000001000000;
		8'd195: 64'b1000000000000000010001000000000010000001100100000000110000100000;
		8'd196: 64'b0000000010000000000000000000010000000100010000000100000100010000;
		8'd197: 64'b0000000000000010000000001010100000000100000000100011000000000000;
		8'd198: 64'b0000000000000000100000100000000001100000010010100000000000011101;
		8'd199: 64'b0001100000000000000000000000000000000000100010000001000001100001;
		8'd200: 64'b0000000100000001000010000000100000000000000000001000000000000000;
		8'd201: 64'b0100001001000000000000001010000000000000000000001010001000000000;
		8'd202: 64'b0000000100000000011000000000100000000000110000011000100000100000;
		8'd203: 64'b0000010010000000000001000100000000000100000000000001000000000000;
		8'd204: 64'b0000000000000000000000000000000010000010100000000001000000001100;
		8'd205: 64'b0000010000000100000100110000000000000000000000000000000010000000;
		8'd206: 64'b0100100010000000101000000000000100010000000000000010010000000000;
		8'd207: 64'b0000110000001000001000000110000000000000100000011000010000000000;
		8'd208: 64'b1000100111000000000000000010000000010000000000000010000000000001;
		8'd209: 64'b0000000010001000000000100000000000000000000000000000000100000000;
		8'd210: 64'b0000000000001001100000000000000000100010000000100000000000000000;
		8'd211: 64'b0000001010001001000000000000000101100100000000000001000000000000;
		8'd212: 64'b0000000000000000100000010100000010100010101000000100000001000000;
		8'd213: 64'b0001001000011000000001000000000000000000001000000010000001000010;
		8'd214: 64'b1000000000000000000000000000000000000000000000100000000000010000;
		8'd215: 64'b0100001100000000000000001000001000100000110000000100100000100000;
		8'd216: 64'b0101010000000010100000000000000000000000000000000000010000000000;
		8'd217: 64'b0000000100000100000000000000000011000000000000100000010000000100;
		8'd218: 64'b0000001010100000000010000001000000000000000110100001010000000100;
		8'd219: 64'b0000100100000000000000000010100000001000000001000000000000010001;
		8'd220: 64'b0000000000000000000000000010000000000000000010000000000000001001;
		8'd221: 64'b0000000000001100000100000100000000010100000000010001000000000001;
		8'd222: 64'b0010100000000000000000100000001100101000000010101111000000000000;
		8'd223: 64'b0000010010000000100000010000000000000110100000010000000000000000;
		8'd224: 64'b0010010000000000000000000010000000000010001000000001001100000010;
		8'd225: 64'b0010001010000000100000000000110000000000000000000000000010000000;
		8'd226: 64'b0100100000010011100000000000000000001000000000000000000100000000;
		8'd227: 64'b0000000000000000010100000000100000001000000000100100001010000000;
		8'd228: 64'b1001000000000000000000101000000000000000110000000000000110000000;
		8'd229: 64'b0000000010100000000000100000000000000000000010000000100000000000;
		8'd230: 64'b0000001000000001010000000000000010000001000001110000000000001000;
		8'd231: 64'b0000000000000100000000101000000101001000000000000000000010000010;
		8'd232: 64'b0000001000000000000000001001100101001000000000001100000000000000;
		8'd233: 64'b1000100000100001000000000000000000000000000010000000000010000000;
		8'd234: 64'b0010101011000000000000000000000000100000000000000100001000000000;
		8'd235: 64'b0000000001000000000000000010010010001000000001000001100000000000;
		8'd236: 64'b0100000100010000000001000000000000001100100100000100000000000010;
		8'd237: 64'b0000000000000000000000000011000010010100000000110100000100001000;
		8'd238: 64'b0010000000010000100010000000010000000001010000010000000010001001;
		8'd239: 64'b0000000000000000100000010000000000000000100000001000001000000000;
		8'd240: 64'b0101000000000000000000100001000000010000000000100000100100001001;
		8'd241: 64'b0000000000001011010000001000100000000000000010010000000000010000;
		8'd242: 64'b0000000110000100000000000000000000100000001000100001010000001000;
		8'd243: 64'b0000001000100010000000000000001000001000000010000110000000000100;
		8'd244: 64'b1100000000001100000110000001000001000000000000010000001000011000;
		8'd245: 64'b0000100000010000000001000100000000000000001001000000000010000000;
		8'd246: 64'b0000100000000001000001000000000000100000000000001001000000000000;
		8'd247: 64'b0000000000000000000000100000000100000000001100000000001000011000;
		8'd248: 64'b0000000000001000000000000000000000000101000000010000001100000000;
		8'd249: 64'b0100000000010001000000000010000000000100100000000100000000000001;
		8'd250: 64'b0100000000000000000000000000000000010000000000000000010000000000;
		8'd251: 64'b0000010001000000100000000000110000000001100001000000000000000000;
		8'd252: 64'b1000000000000000110010000000100000000001000100001011000000100000;
		8'd253: 64'b1000000000000000000000000001110000000010010000000000001100000100;
		8'd254: 64'b1000000000011001100001000000000010000000001000100001010000000110;
		8'd255: 64'b0000000000000000001000010000000000000000000000001000100000010000;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page1(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1000000001001000001111000110000000000000000101000001000001100001;
		8'd1: 64'b0001001010000010000001100000100101000100101001010010000010001101;
		8'd2: 64'b1010100100000000000010000001001000110100100000100000011110000011;
		8'd3: 64'b0001001000010000111000000001000010010000000100000010000000010010;
		8'd4: 64'b0110000000000100000000000110100001100000100001000000001000101100;
		8'd5: 64'b0000000000100000110000110100000001111100000001001101001101000100;
		8'd6: 64'b0001100001000000000000110000000001001000010010100010101100100000;
		8'd7: 64'b0000000101000001010000000000100000101100000010000000000100000000;
		8'd8: 64'b0000010000011000001100000001000000101001000111000011101100001000;
		8'd9: 64'b0100100010000000000001010000001010001000000000100000001100010100;
		8'd10: 64'b0000000001001000010100100011101000000000011100001000000011110000;
		8'd11: 64'b0000000011000000010000000100001000001100000010000110110100100110;
		8'd12: 64'b0000010011110010100010100000011101001010010111001000100000100101;
		8'd13: 64'b1011100001000010000011000000000000010000000000000000101001000001;
		8'd14: 64'b0000001100000000000010000100010000000000010100100001010000001100;
		8'd15: 64'b0010010010000000001010000000000000010100000110010000010001100010;
		8'd16: 64'b1100000010000000100000010000000001000000000000101000010001010000;
		8'd17: 64'b0001001100000100000000000000000000000001000001001100000000000001;
		8'd18: 64'b0000100000000110000000110000000001010011000100000000001000000000;
		8'd19: 64'b0001100000000001001000001001001010000000011010011100001000000100;
		8'd20: 64'b1010000000011000000100000110001100000000101011001000100000100000;
		8'd21: 64'b0000000001000010101000010110000010000000000000001010110010001101;
		8'd22: 64'b0000000000000010010001001000101010000100000111001000100010000011;
		8'd23: 64'b0000000000001000110000000111100000100000001000011100001101010111;
		8'd24: 64'b0000101000000100100000011000000100100000001010000010011010100000;
		8'd25: 64'b0001000000000000000011011011010001100010000001010001001010000010;
		8'd26: 64'b0101000001000101100000001000010000001010101010000000001000000000;
		8'd27: 64'b0100000101000110010001000101010001001000111100000110000101000100;
		8'd28: 64'b0000101000000100000001000001010001110010101000000000010010000100;
		8'd29: 64'b0001100111010010000001010000010100001000000000000000110000101000;
		8'd30: 64'b0001010100000010000000010001000001100000000001000000000010000000;
		8'd31: 64'b0000000100000100000001011001000000110000000000000000001000000011;
		8'd32: 64'b0101100100001000000000001100000000111011110001110000000001010000;
		8'd33: 64'b0001000000010101001001010000000001101100000001011000100000000100;
		8'd34: 64'b0000100100000011000001111000000001000011000001000000001100000000;
		8'd35: 64'b0000010100000011000000000010000111000011100000000000001100001100;
		8'd36: 64'b1000000000000000101000101000110000000011000000000010000000000100;
		8'd37: 64'b0100100000000000000000000100000010010000101000000011010110100000;
		8'd38: 64'b1011110000001000000001000100001001000010000000011000010100000010;
		8'd39: 64'b0011000010001000000100000000010100010101010011001100001000001001;
		8'd40: 64'b0101001100000000000000101010100100111010000000000010010010010111;
		8'd41: 64'b1001100100000010000000000001000000001010100001000000101000000000;
		8'd42: 64'b0000001001001100010000010000001010000000000010000100011000001001;
		8'd43: 64'b1001010000000100101000100000010000011001001000100001000000100100;
		8'd44: 64'b0100001000000000000000110000001111000000010010000000000010010010;
		8'd45: 64'b0111100000010110110101010000000101010001010000100001000000100010;
		8'd46: 64'b1000000000101000001000011101011000000100001010001000001001001000;
		8'd47: 64'b0100010001000000000000000010000100110100000000000010000000001000;
		8'd48: 64'b0000011001101000101000000100000000001000000100010010100000001101;
		8'd49: 64'b0110000000000000000010110010000100001000000000011000100000010000;
		8'd50: 64'b0001001000011000010100000010000100100110110011010000100000001011;
		8'd51: 64'b0100110100000000001000000110000001000000000000010000100110101000;
		8'd52: 64'b0000010001000001100101100000000100001001001001010100000001010001;
		8'd53: 64'b0001100010000001001101000100000001000000001000010000100101100110;
		8'd54: 64'b0000010110110000010000000110001000100110000000100000000000111000;
		8'd55: 64'b0000010011000000010000000001001100001000000110110000001101110101;
		8'd56: 64'b1100001001000000001011000000000000000000001001010010000010001000;
		8'd57: 64'b0000000010001100000000100000000000011010011000001110000100000000;
		8'd58: 64'b0000000011100000010100000100000000000100010000000100100000100110;
		8'd59: 64'b0010001000010000000000010100000000100010010001000011010100010010;
		8'd60: 64'b1010001000000111011100000111011100010000000010000001001001001000;
		8'd61: 64'b0100100000000000010000000011000110101110001000000000010000010100;
		8'd62: 64'b0100001000001000100100010101000100000010001001001001000001010100;
		8'd63: 64'b0011000000001000000100000000110101000010000000000000000101000001;
		8'd64: 64'b0010010000100000001000100001001010100000100000010000001110100000;
		8'd65: 64'b0010000000000100111000000011100000000000000000000100000010000100;
		8'd66: 64'b0110000011000010000110000101000100000000010010010010000011000101;
		8'd67: 64'b0000111000110001000011100000110000010010000000000000001000011000;
		8'd68: 64'b0000010000000100000001001000001000000000110010011000010000000000;
		8'd69: 64'b0101000000000001000000000001101000001100001000111001000000000000;
		8'd70: 64'b1000010010010000000000001000000000000000010100010000000000110110;
		8'd71: 64'b0010000000000110000000000000101000000100001001000000010000001100;
		8'd72: 64'b0000001000000010100000001000000000001010101000011000001000000100;
		8'd73: 64'b1100000010000000000000001100010101010000010010100001001001000011;
		8'd74: 64'b0000001011000001000010000000001110010110000100000100100010010100;
		8'd75: 64'b0000000101001001000010000001100000000000000110000000100001001001;
		8'd76: 64'b1000100011010100000000000001000001000000100101001000010000110010;
		8'd77: 64'b0001000010010011010000010110001010111100100100100000100110000110;
		8'd78: 64'b0100100000001000110000000101010000001100100011001101010000001101;
		8'd79: 64'b1000010010100000110010000000000100000000000010110010000000000000;
		8'd80: 64'b0011000000010100000001000001010000000100000101000010010100000010;
		8'd81: 64'b1000000010111000010000010000100001000101010000000010000000000001;
		8'd82: 64'b1100000000100000000000001001001000010011100000000000010000000000;
		8'd83: 64'b0000001010000011111010010000000000011000100000001000000100100110;
		8'd84: 64'b0100000010101001101110010000000100000001011100000100000010001100;
		8'd85: 64'b0000000000000100000000000010010000100010111101000010111101100000;
		8'd86: 64'b0010010000000100001101100100010000101101010000011011110100001100;
		8'd87: 64'b1001100000000000100001011010000000001000011011000010000000001000;
		8'd88: 64'b1000000000001010110010010000011000100000101001100000100000001100;
		8'd89: 64'b0100000000010000010100000101000000001100110000001010000000100000;
		8'd90: 64'b1001010010110110000000000001000010010011001100000010001101010100;
		8'd91: 64'b0000010000100001010000000001000000110010100000000000000000000010;
		8'd92: 64'b0011000111100010001000000000000000111001000000000010000000000001;
		8'd93: 64'b1010110000000000100000000010000000001101001000000000001001000010;
		8'd94: 64'b0101000001011010000110010001100000010001001100000000101000000010;
		8'd95: 64'b1101000110000001000000000010010000010100001010000000010000010011;
		8'd96: 64'b0010001100010010000000001000001000011000110111000001010110010010;
		8'd97: 64'b0000111000011011000000100000001001101100001000000001000000000001;
		8'd98: 64'b0000000000101000000000010110000001000000001000010100010001001001;
		8'd99: 64'b1001001000000000110010000100011000000100100001000100001100000010;
		8'd100: 64'b0000100100001000100010000000101000010000000000000101010010000001;
		8'd101: 64'b0010000010000100001011000100000001010000001001010010001000000000;
		8'd102: 64'b0011001000011000000100100000010001100010000110100001000010000000;
		8'd103: 64'b1100000000000000001110100000000010001000000000000100010101010000;
		8'd104: 64'b0000011000000011000101010000000010100000101000100100001110011000;
		8'd105: 64'b1001000000000000010010111110100011100110100100010101100100000000;
		8'd106: 64'b0100101100010001010000100100001000010010001000000100001100001000;
		8'd107: 64'b0100000100010011000010100000100001011000000001000100000000011000;
		8'd108: 64'b1000100001000000001001000010100011010000001101100000010000001010;
		8'd109: 64'b0010010000000000000010010010011000010000001010000100000100000110;
		8'd110: 64'b0001000010001011000100000010111000001000101100101000000001100000;
		8'd111: 64'b0101101010000000000010010000011000100001100100110011000100110011;
		8'd112: 64'b0001001000010100100001000000010001010110001100000010110000000011;
		8'd113: 64'b1001000000001001000100001100000001010000000001110000000000010010;
		8'd114: 64'b1001100010000000000000001001100100101001000010000000010100010001;
		8'd115: 64'b0100000110001000010100010000000001100001001100100001000000000010;
		8'd116: 64'b0100000000100101000010010000000000000001000100100010110000101100;
		8'd117: 64'b0000000101110101001010100110000001000000010011000000110100000101;
		8'd118: 64'b0110001000000001000000001000100000010000101000010000001000100110;
		8'd119: 64'b0100111000010010000001010000001010000110100110101000011110010010;
		8'd120: 64'b0000000000110011011000000001010000100011101000000100010000000001;
		8'd121: 64'b0011001011000100010000100000100001000000010000000000000100000000;
		8'd122: 64'b0010000000000100001101000000100000100000010000010000000001000100;
		8'd123: 64'b0100000010100000000110001000000000100000010010010010000000100010;
		8'd124: 64'b0000100000010010100001001010000000000000001000000000000101011010;
		8'd125: 64'b0111000000011000000001000001010000101000111001000010010000100010;
		8'd126: 64'b0010000000111010000000000000001001000000100010001010000110000101;
		8'd127: 64'b0000010000000110011010110100010100000001001000000000000000000001;
		8'd128: 64'b0000110010110100100011000100001100010000000001001100110000010010;
		8'd129: 64'b1000000110010010110100000101000001011001001000000010000101000000;
		8'd130: 64'b0000000100001000000100000001100110001011001000000001011000011100;
		8'd131: 64'b1101000011000000001110000000000010001011000000011000111000100000;
		8'd132: 64'b0011010010101000100010011011000100010001100000001111010100000001;
		8'd133: 64'b1001101000100000001010100101100000011001000110000000000000000000;
		8'd134: 64'b0000100011001000010000100110000000100001101000100100011001000000;
		8'd135: 64'b0010000000100000000000100011000000100000000000010110000000000000;
		8'd136: 64'b0010000010000000100000001010000001000000100010000010010010000010;
		8'd137: 64'b1000011111000000101001010011001000010000000101000000000100100001;
		8'd138: 64'b0101000101010101001100100000110001001100010001110100000001001100;
		8'd139: 64'b0001010010110001001010100111100010000000001010000110100000000100;
		8'd140: 64'b0000000000001000000010011000000100000000100000100000101000011000;
		8'd141: 64'b0000000000100000000010011000001010010000001100000010011110100001;
		8'd142: 64'b1100101000111010000000000001101011101000000101100000100000010001;
		8'd143: 64'b1110100011000000000000001110001100001000001000110000000001000101;
		8'd144: 64'b1000000101101100000000011101100010010001000001010000000000010000;
		8'd145: 64'b0011100010010101000001000101010100000110000000000100001101110110;
		8'd146: 64'b0100010001000110011000000100000000101010000101100000000111000101;
		8'd147: 64'b0110000000000100100000001000001100100011100000011100000010000000;
		8'd148: 64'b1000011000000001010100010000000000001000001000000000101000000100;
		8'd149: 64'b0010100001000010000000011111011000001000001000000000000001000010;
		8'd150: 64'b1010100010000100100000000011001100100000010100000000010010100000;
		8'd151: 64'b0100000000010011100111000000100010000100000000000011000101000000;
		8'd152: 64'b0000100000000001101010100110001010101110000111100000001000001010;
		8'd153: 64'b1101011010010000100100011000000000011000101000000001010000110001;
		8'd154: 64'b0000010100000000001010001111000000000100000001001010110000001110;
		8'd155: 64'b0000100000100010010101000000000000010000000001010100000000010000;
		8'd156: 64'b0000000101011001100000010001000000001000000001100011000000011010;
		8'd157: 64'b0111000100001000110100000111000011010000000000000001000011100000;
		8'd158: 64'b0100100000000101000001001000000001100000000010000000000000110010;
		8'd159: 64'b1000110101000000000100101010000000100000001000000010010001000010;
		8'd160: 64'b0000110000000010000000010011000000000000110001000000000000001000;
		8'd161: 64'b0000000000010010100000001010100010101100000000100000000000101000;
		8'd162: 64'b0110011011001000010101001100000000100010010000000100100101100000;
		8'd163: 64'b1111010001010010100001001110101001000000000100010000010000101000;
		8'd164: 64'b1000000000000001000100010000111100000001000000010011000110001000;
		8'd165: 64'b0000111000000101100010100001001100101111010011010000000000001001;
		8'd166: 64'b0000010000000001000001010001111001010001101001010011001100100000;
		8'd167: 64'b1010010010000000001000101000001111100000000000000000100001000000;
		8'd168: 64'b0001001000001000110101000000100010110100000000000001000001001100;
		8'd169: 64'b0100011010000000010100000000000110000000100000001100100010000101;
		8'd170: 64'b0000001000001100001000001110001100000000010010000000000101000000;
		8'd171: 64'b0011100011000100000000001010011100000110010010000000000000000000;
		8'd172: 64'b0010100000101111001010011101000000101001000010110010000001010000;
		8'd173: 64'b0001010001000000000000000100001001000001110000001000000010000010;
		8'd174: 64'b0000000101100000100101000010010000110000100011010100110000011000;
		8'd175: 64'b1011000010011000001000000000001010010000000110011010100010000010;
		8'd176: 64'b0011000100011101011010000100001101010101100000000011000000101010;
		8'd177: 64'b0010100010000000100001000001100000010000000001001000100011010100;
		8'd178: 64'b0010001110000000001000000000100010000000000000000000000100000001;
		8'd179: 64'b0010010010000100011000001001001101011001101000100010001001110110;
		8'd180: 64'b0010001000000000000000010000000010000000000010000000010000000010;
		8'd181: 64'b1001000110010000001000001100000010000001001000100010000010000000;
		8'd182: 64'b0000000011111000010010101000000000101011011100100000000000000000;
		8'd183: 64'b0011000010000000000010000000000000001001101111001100000110001100;
		8'd184: 64'b0110000100100000001001001000000101001010000001000000000010000000;
		8'd185: 64'b0001000100010001011000000000001001001100010101000001000100000100;
		8'd186: 64'b0000001101100010000010001001001010001000000100000100000101001001;
		8'd187: 64'b1001000101100010000010000000000011001100000000010001011010000110;
		8'd188: 64'b0010001000001000000011001001000000000100010010100001001000000000;
		8'd189: 64'b0100000000010011100000000000010000000000000000001000000000101110;
		8'd190: 64'b0000000100010000010000010110000001000100001101100001010001000001;
		8'd191: 64'b0100000001101000101001100001000100010010010000100001101000000000;
		8'd192: 64'b0110011001000101001000100010101001000110000000110101010000100000;
		8'd193: 64'b0101000001100101010000101000110000001110000000100001000000000001;
		8'd194: 64'b1001000000000101010100000010000011010111100001010001000001001000;
		8'd195: 64'b1000000000000000110001000001100010000001100100000000110000110100;
		8'd196: 64'b0000000010000001000000000000010000000110010000100101000100011000;
		8'd197: 64'b0001001000000010000001001010100000000100001101100011001000100001;
		8'd198: 64'b0000000000000000110001100000000001100001010010101100010000011101;
		8'd199: 64'b0101100011001000000000000000000100010010100010000101000001100001;
		8'd200: 64'b0001000110010001000110000010100000000000000100101001000010000100;
		8'd201: 64'b0100001001000000000000001011000000000000000000101110011000000000;
		8'd202: 64'b0000000100101010011000010010100000000000110000011000100000110010;
		8'd203: 64'b0100010010000010000001010100010001000110000000100001000001100000;
		8'd204: 64'b1000000000100000100000100000000010001110100000001001000010001100;
		8'd205: 64'b0000010000000100000100110000000000000000010000010000000010000100;
		8'd206: 64'b0100100010000001111001000000000100010000000000000010110000100000;
		8'd207: 64'b0000111000001010001100000110000000000100100000111010011101000000;
		8'd208: 64'b1001100111001001001100000010000000010001000000011010010000000001;
		8'd209: 64'b0001000010001010000010100100000011000000010000000000000100000000;
		8'd210: 64'b0010000000011101100010010001100000100010000100100000100001001000;
		8'd211: 64'b0100001010001001000100000010100111111100000100000001000010111100;
		8'd212: 64'b0000011000000000110101011100001010100110101000010100000001000000;
		8'd213: 64'b0001001000011011000001010000001000000000001101101010100001011010;
		8'd214: 64'b1000000100000000001010000000000000100100000000110000000000010000;
		8'd215: 64'b0110101111000000000000001000001000100000111000010100100000100010;
		8'd216: 64'b1111010000001010100000000101001010010000000000000000010001010110;
		8'd217: 64'b0000000100000100010101000001000011000000000000101000010000000100;
		8'd218: 64'b0000001010110010000011000011010000000000000111111001010000000100;
		8'd219: 64'b0001100100011000000000000011100000001000100011000000000000010001;
		8'd220: 64'b1001000000010000000000100011010000000000000011000010100000001001;
		8'd221: 64'b1000000010001100000100000100000010010100000010010001000000000001;
		8'd222: 64'b0010101000101000000001100000101100101010010010101111000001000000;
		8'd223: 64'b0000011010010000100000010000000000000111100000010000000010000000;
		8'd224: 64'b0010010010100000001101101010000000000010001000000011101110000010;
		8'd225: 64'b0010011010000000100100100000110010100000000000100000001010000000;
		8'd226: 64'b0100101000010011100000000000000101001000000100100100000100000000;
		8'd227: 64'b0000110000000010010101000000101000001000000100100100001010100000;
		8'd228: 64'b1001101110001000000000111000001000000001110110000010000110001000;
		8'd229: 64'b0001000010100100000111100000000000000000000010001000101000010000;
		8'd230: 64'b0001001001001001010000000001001010000011000001110000000010001000;
		8'd231: 64'b0100100000000100000010101000000101001000001000100000101010100010;
		8'd232: 64'b0010001000000000000001001001100101001010000001101100000010100100;
		8'd233: 64'b1000110000101001100000000010000010001010011011000000001010100000;
		8'd234: 64'b0011101011000000010000000001000000100011000000010100101000000010;
		8'd235: 64'b0100100001000000110100000011010010001011010001000001100000100000;
		8'd236: 64'b0100000100010000010001000010000010101101101100000100000000010011;
		8'd237: 64'b0100100001100000000000001011001011010100000011110100000100001000;
		8'd238: 64'b0010010010011000100110000100010000001001010000010110000010001001;
		8'd239: 64'b1000100000000000100110110000000010000000100000011000011101100000;
		8'd240: 64'b0101000000000000010000100001000010010000010000110000100100001001;
		8'd241: 64'b0000000001001011110000101000100000000000000010110100000000010100;
		8'd242: 64'b0000000110000111010000000000000000100000001001100001010010011010;
		8'd243: 64'b0001011001100010010000100010001100111001000010000110001000100111;
		8'd244: 64'b1100000000001101000110000101000001000011000001010010001001011000;
		8'd245: 64'b0000100000010000000001000100000010000000001111000000000010000100;
		8'd246: 64'b1000100000000001010101001000001000100000000000001001000100000000;
		8'd247: 64'b0000000000100000000001100000010100001100101101000100001000011000;
		8'd248: 64'b0000011000001010001000000001011100000111000000010010001101000000;
		8'd249: 64'b0100000000110011000000000011000000000100101100000100000000010001;
		8'd250: 64'b0100100000000010000001000000101000010100100000000000010000000000;
		8'd251: 64'b0000010001100011100100000000110001000001110001000000010000000100;
		8'd252: 64'b1000000100000010110010000010100000101001000100001011000000100001;
		8'd253: 64'b1000101100001010100000000001110101000011010111000010001100000101;
		8'd254: 64'b1000110010011001100001001110000110110000001000101001011001000110;
		8'd255: 64'b0000000000001000111000011000000000100010000000001000100000010010;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page2(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1000010001011000101111100110000100000000101101001011000001100011;
		8'd1: 64'b0001011010100110110001100010100101100100101001010110001010101101;
		8'd2: 64'b1110110110000000000010100001001100110100100100100000011110010111;
		8'd3: 64'b0001001000010000111101000011000010010100000100000010010000010010;
		8'd4: 64'b1110000001100100010000010110100001100000110001000010011000101100;
		8'd5: 64'b0001000010100000110001110101010001111101000001011101001111000100;
		8'd6: 64'b1001100001100000000000110001000001001000011010101110101100101000;
		8'd7: 64'b0000011101000001010010000000100000101110000010100000000100000000;
		8'd8: 64'b1001111010011101001100000001000000101001001111100011101100001000;
		8'd9: 64'b1110100010000000000011010000101010001011000010101010001100010100;
		8'd10: 64'b0100001001011010010100100111101000000010011110001010000011111000;
		8'd11: 64'b0010100011010000010000001100001100001100001010100110110100111111;
		8'd12: 64'b0100110011110010100010100010011101001010010111001001101000100111;
		8'd13: 64'b1011100001000010010111000100010000011000000100000000101001000001;
		8'd14: 64'b0001001100110010000110110100011001000000110100100011010000111101;
		8'd15: 64'b1111010010000000001010000000000000010110000111010000110001100011;
		8'd16: 64'b1100000010011000100000010100000111000000100010101010010001010001;
		8'd17: 64'b0001001100001100010010000100000100100001000001001100000010000001;
		8'd18: 64'b0100111010000111000110110100101001010011000100100000101100001000;
		8'd19: 64'b0001100100010011011000011001001010010001011011011100001000011100;
		8'd20: 64'b1010000000111000001110000110101110001000101011001011101000101000;
		8'd21: 64'b0000101011100010101000111110001010000010100000101010111011001101;
		8'd22: 64'b1000000000010010010011001010101011000100010111101000100010001011;
		8'd23: 64'b0010000000001001110010000111100101100001101100011100101101010111;
		8'd24: 64'b0000101000001100100000011000000101101000101110001110111010100111;
		8'd25: 64'b0111000000000001000011111011010001100010000001010001001010000010;
		8'd26: 64'b0101010001000101100000101000010010001010101010000000101111001000;
		8'd27: 64'b1100101101011110010001010101011011001011111101000110100101011100;
		8'd28: 64'b0000101000100100001001111111010001110010101001100000110011001100;
		8'd29: 64'b1001100111010011100011010010011110001111100000000000111000101000;
		8'd30: 64'b0001010100000010010000010101001001100000010001100000001010000000;
		8'd31: 64'b0000000100010100000001011101100001110000000010000100001000101011;
		8'd32: 64'b0101111110101010000000001100100010111011110001111100000001010100;
		8'd33: 64'b0011001001011111101111010000001101101110000101011010100000100100;
		8'd34: 64'b0100100110000111000001111110011001100011100001000000011100100010;
		8'd35: 64'b0000010101000011010000010010000111000111110010010001001100101100;
		8'd36: 64'b1100010000000000101000111000110100011011010011000011000011000101;
		8'd37: 64'b0100100000000000001010001110000010010000101000000011010110110000;
		8'd38: 64'b1111110000111000100001010100001001001110010000011001010100000011;
		8'd39: 64'b0011001010111100100100000000010110110111110011101100001100001001;
		8'd40: 64'b0101001100000001000001101010100101111010000000100010011010010111;
		8'd41: 64'b1001100100010110000010000001100000001010110001001000101100001000;
		8'd42: 64'b1000001011011100011110111000001010101000011010000110011100001001;
		8'd43: 64'b1001010100001100111000100000010010011101001001101001010000100100;
		8'd44: 64'b0100001000000001000010110001001111000000010010001001000010011011;
		8'd45: 64'b0111100100010110110101010000001101110011010001110101100000101010;
		8'd46: 64'b1000000000101001001000011101111110000100001110001000001101001100;
		8'd47: 64'b0100010001010000000000100010000101110101000011000010001000001000;
		8'd48: 64'b1000011111101000101000000100010100101000010100010010100100001101;
		8'd49: 64'b0111000001000001000110111110000100011010010000011000101000010000;
		8'd50: 64'b0001101001011001110110010010110111110110110011010000111010001011;
		8'd51: 64'b1110110100000000101001100111000101000001110000010110110110101000;
		8'd52: 64'b1001010001000001100101100000000101011001001001010100000001010001;
		8'd53: 64'b1011100011000101001111000100000001110000001001110001100111101111;
		8'd54: 64'b0000011110110100011001100111001000100110000101100000010001111100;
		8'd55: 64'b0000110011100110010000010001001110011000000110110000001101110101;
		8'd56: 64'b1100001001001000101011000000000000000010001001010010010010001000;
		8'd57: 64'b0001000010011101000000100000000001011010011010001110000100000001;
		8'd58: 64'b1000000111100000110100001100001010010100010000000101100000100110;
		8'd59: 64'b0010011000011001000000010100000001100110011101010011010100110010;
		8'd60: 64'b1010011000100111011100100111111100011100011010000001101001001011;
		8'd61: 64'b0110100000110000011000000011000111111110111010100010010010010100;
		8'd62: 64'b1100011010001000101100010101100101100010111001011001000101010111;
		8'd63: 64'b0011000010001100000100001000110101000010000100000000100101001001;
		8'd64: 64'b1010011000100010001000110001001010100000110000010000001111100011;
		8'd65: 64'b0011100010000100111000000011100000010010100101000101000011011100;
		8'd66: 64'b1110001011001010001110000101011110110000110011010010000011000101;
		8'd67: 64'b0000111000110001000011111000110000010010010100000000001000011000;
		8'd68: 64'b1000010001100101001001001000001010000000110010111100010110001000;
		8'd69: 64'b1101100000000001100000000011101000001101101000111001000000000010;
		8'd70: 64'b1000110110010000000010101001001000011000010100011000100000111110;
		8'd71: 64'b0010000111000110000000010000111000100100011011000000011010001110;
		8'd72: 64'b0000001111001011101100001001000000001010101001011000001110000100;
		8'd73: 64'b1110001010000000000110001100010101110011111010100001101001000011;
		8'd74: 64'b0001001011010011010010101110001110111110011100000101111010010101;
		8'd75: 64'b0100100101001001000010110001100000100001000110001000100001001001;
		8'd76: 64'b1000100011010100000101001001000001000100100101011000010010110110;
		8'd77: 64'b0001000010010011010000010110111011111100110100101100100111000110;
		8'd78: 64'b0101100100011000110010000101110010001100100011001111110000001101;
		8'd79: 64'b1000011010100001111010100001001100000100000010110011010000000001;
		8'd80: 64'b0011010110110100000101000001011010110101000101100010010100100010;
		8'd81: 64'b1000000111111011010001010000100101000101011000000110010000001101;
		8'd82: 64'b1110000000100000111011001001001000010011100000000001010000010000;
		8'd83: 64'b1000001110000111111010010000000010011000101010101110000100101110;
		8'd84: 64'b0100000110101111101110110000110101000001011101000100100010001100;
		8'd85: 64'b0000110000100111000000000010011000101010111101000010111111100000;
		8'd86: 64'b0010010000001100001101100100010100101101010001011011110100001101;
		8'd87: 64'b1111100000100000110001011010000100101000011011000010000000001010;
		8'd88: 64'b1000000111101010111010010001111000100000101001100110111000001110;
		8'd89: 64'b0100010000110000110100010101010000001100111000001010010000100000;
		8'd90: 64'b1001010110110110000010010001100110010011001110000010001101010100;
		8'd91: 64'b0001010100100001010000000001001010111110100000000000000000000110;
		8'd92: 64'b0011010111100011111000001101000100111001000000001011100010000001;
		8'd93: 64'b1010110010001000100000001010100010101101001000000001001001001011;
		8'd94: 64'b0101001011011010100111110011100001011101101100100000101000000010;
		8'd95: 64'b1111010110000011000001010010010000010100101010000000010000010011;
		8'd96: 64'b1011101101011010100101011001001000111001110111000001011110010010;
		8'd97: 64'b1000111000111111100100100000001001101111001001000001110000000001;
		8'd98: 64'b0100000001101001010100110110010001100000011000110100111001101011;
		8'd99: 64'b1001001001010000110010100110111000000100101101000100001101010010;
		8'd100: 64'b0000101100001000100111001010111000011000100000000101110010000101;
		8'd101: 64'b1010110010011111011111001100010101010000001001011011011010001000;
		8'd102: 64'b0011001000011100000100100000010001101010010111100011001010001000;
		8'd103: 64'b1110000011010000001110100001000010001100000100000100011101010000;
		8'd104: 64'b1100011000000011000111110000000010100000101001100100001110011000;
		8'd105: 64'b1111101000101000010010111110100011100110100110010101100100000100;
		8'd106: 64'b0100101101010001010001100100101001111010011000000100001100011010;
		8'd107: 64'b0100010100010111010010100000110011011100000001000110000101011000;
		8'd108: 64'b1000101011000100001001101010100011010010001101100000010000001010;
		8'd109: 64'b1110010100001000010010010010011000010010001010000100100110000110;
		8'd110: 64'b0001010010101011000100000011111010001000111100101001001001100000;
		8'd111: 64'b0101101010000100000010010000011000110001100100111011100100110011;
		8'd112: 64'b0001001000010101100111100000010111010110001110000010110000000011;
		8'd113: 64'b1001000000001011000100001101001001010100000011110000000001010011;
		8'd114: 64'b1011110010001000000000001001100100101011000011000001110110010001;
		8'd115: 64'b0100000110111001010100010000000001110001001100100011000000100010;
		8'd116: 64'b0110000000101101001010010000000000110011000100100011110000101100;
		8'd117: 64'b0000011111110101001010100111000001000100010011100000110111010101;
		8'd118: 64'b0110101000000001010000001000100000010010101010010000001110101110;
		8'd119: 64'b0100111000010110000101110001001011101110100110111000011110010010;
		8'd120: 64'b0000000000110111011000101001011100100011101101010100111000100011;
		8'd121: 64'b0111101011010100110010100110101011000100010000000110001100100000;
		8'd122: 64'b0010001000100101011101000000111000100010011000010000001001000110;
		8'd123: 64'b0100000010100000010110001110100000100000010010111110000001100110;
		8'd124: 64'b0001100000110010100001011011100001000001101000100000000111011010;
		8'd125: 64'b0111100000011000000101000001010100101000111101100010010000100011;
		8'd126: 64'b1010001100111010000101000000101011000011100010001110100110000111;
		8'd127: 64'b0001010101000110111010110110010100000101001000000000000100100101;
		8'd128: 64'b0000110010110110100011000100001100111000010001001100111000010011;
		8'd129: 64'b1001000110011010110111010111000101011001001000010010001101000000;
		8'd130: 64'b0100000100111000100100000001100110011111111001001001011000011101;
		8'd131: 64'b1101100111010001101110001010000010001011110000111001111000100000;
		8'd132: 64'b0111110011111110101010011011000100010001100000101111010110000111;
		8'd133: 64'b1001111100110100001010101101100111011011000110010100011001000000;
		8'd134: 64'b0000110011001000010001100111000011100001101010100110111101000000;
		8'd135: 64'b0111011000110010000000100011100000100001111000110110100010001000;
		8'd136: 64'b0010000011000000100000011110000001101000110010010010010011000110;
		8'd137: 64'b1101011111010000101001111011011000010000110101010001000100100101;
		8'd138: 64'b0101010101010101111100101000110011101100010001110110000001001100;
		8'd139: 64'b0101010010111001101010100111100010000100001010000110100101100110;
		8'd140: 64'b0000101010001100100011011000000101000000100001100000101011011000;
		8'd141: 64'b0100000110111100000110111000111010010000001100000010111110100101;
		8'd142: 64'b1100111100111010011110000011101111101010000111100010101001110001;
		8'd143: 64'b1110100111000000000100011110001100011000001010110000001001000111;
		8'd144: 64'b1000010101111101100000011111100010010101100101011001011000010100;
		8'd145: 64'b0011100010010101010001010101110100000110001000000100001101111110;
		8'd146: 64'b0110110011000110011000000110100010101010000101100000100111010101;
		8'd147: 64'b0110100000000100100000101010001110100011101000011101000010000000;
		8'd148: 64'b1000011010000101010100010001100000001000001000000001101000000100;
		8'd149: 64'b0010100001100010000000111111011000011001001001000000101001000110;
		8'd150: 64'b1110100010010100101001000011001110101000010101000000111110110000;
		8'd151: 64'b1100000100110011100111000100100010000100000000001011010101000000;
		8'd152: 64'b0010101000000101111010100111011110111110000111111000011001101111;
		8'd153: 64'b1111011110010001100100111001011011011000101100010001011010110001;
		8'd154: 64'b0110010100000000011010001111001001001101000001001010111101001110;
		8'd155: 64'b0000100100100010110101010000100001011000000001010100110000010000;
		8'd156: 64'b0100000101011101101000110001001000001000010001100111111100011010;
		8'd157: 64'b0111010110001000110100000111000011010010110000000101000111100000;
		8'd158: 64'b0100100101001111000001001010001101100100000010001100000001110010;
		8'd159: 64'b1000110101100100101100101111000010100000001011100010010111001010;
		8'd160: 64'b0100110000010110100000011111000100000101110001000100000101001101;
		8'd161: 64'b0000000000110010111001101011100010101101000000101000010000111000;
		8'd162: 64'b0110011011011000011111011101001000100110010010000100100111100001;
		8'd163: 64'b1111010001111010100001001111101001000001110100010001010010101000;
		8'd164: 64'b1000100100010001000110010010111100000001000000010011000110001100;
		8'd165: 64'b0101111001000101100011101001001100101111110011010100110110001001;
		8'd166: 64'b0000010000011101000001011011111001010101101101011011111111110010;
		8'd167: 64'b1010010010100001101000101100001111101100000000011000100001001010;
		8'd168: 64'b0011101000101000110101001000110110110110001010000001100001001100;
		8'd169: 64'b0100011110001011010110011000000110010100100010001100100110000111;
		8'd170: 64'b0000101100001110001110101110101100000010010011100000000101001000;
		8'd171: 64'b0111110111101100000011101010011101001110011011010000010000000000;
		8'd172: 64'b0010111010101111001010011111000000101001110011110010000001010001;
		8'd173: 64'b0001011111000001000000010100101001000101110000101100000110000010;
		8'd174: 64'b1010000101100110100111000010010000111100100011010101110010011000;
		8'd175: 64'b1011001010011001001010101101101010010000011110111011100010101010;
		8'd176: 64'b0111010100011101011111001101101101010101100101000011100010101011;
		8'd177: 64'b0010100010010011101001000101100000011000000001001011100011010100;
		8'd178: 64'b0010101111000010101001000000100010000000000000100001010100000001;
		8'd179: 64'b1110110010000100111001101011001101111111101000101010011001110110;
		8'd180: 64'b0010001000000010101100010000000010010010000011000000010001100011;
		8'd181: 64'b1001000110010010001110001100001010011001001010100110000010010000;
		8'd182: 64'b1000000011111000010010111001001000101011111100100000100110001000;
		8'd183: 64'b0111000010001000000110000000000000011001111111001100010110001100;
		8'd184: 64'b0110100100100010001101001000010101001011000001000000000011000000;
		8'd185: 64'b1001010100010001011000000000101001001100010101000001100111000101;
		8'd186: 64'b1001001101100110000010001101101111011000000100000100000101001011;
		8'd187: 64'b1001000101101010001011010000000011001100001000010001111010001110;
		8'd188: 64'b0010001000001000010011011101100000001100110010100001101000000000;
		8'd189: 64'b0110000000010011100000000100010001100000010100101100000100101110;
		8'd190: 64'b0001010110110000010100010110010011001100001111101111011001100001;
		8'd191: 64'b0100000001111000111001100001000100110010010010101001101100110011;
		8'd192: 64'b1110011001001101111000111110101001000111010010110101010001100000;
		8'd193: 64'b0101010001100101010001101000111000001110000010100001110001000011;
		8'd194: 64'b1001001100100101010100000110000011010111100101010101001101001101;
		8'd195: 64'b1000000000010111110001000001110010000001100100001001110000110100;
		8'd196: 64'b0100000010010001010100000000110001000110110110100101000100111000;
		8'd197: 64'b0011011000100010000101001011100011100100001101100011101000101011;
		8'd198: 64'b0000001000101111110001100000000101100001110011101101010000111101;
		8'd199: 64'b0101111111001001010000000110100100010110110010100101010101100011;
		8'd200: 64'b0101001110010001100110010011100000011100010100101101010010000110;
		8'd201: 64'b1101001001010000111000001011000110010000000000101111011000000000;
		8'd202: 64'b1010100100101110011000110010100000101000111100011110100000110010;
		8'd203: 64'b0100011010001010000001010100011001000111000001100011011111111000;
		8'd204: 64'b1011000010100000100100110000000011101110100000001001001010001100;
		8'd205: 64'b0100011000100100000110110000000100001100011000110000000010000100;
		8'd206: 64'b0101100010000001111001001001010101011000100000010110110000100000;
		8'd207: 64'b0010111000001011101101110110001000100100100010111010011101001010;
		8'd208: 64'b1001101111001001001100100010001110110001000000011010010001000001;
		8'd209: 64'b1001000010111010000010110100010011000000010000000000000100010101;
		8'd210: 64'b1010000000011101110011010101111111100010000111101000100011001000;
		8'd211: 64'b0100011010001101100110101010110111111110000100100001110010111101;
		8'd212: 64'b0000011000000000110101011110011010100110101000110100001001000101;
		8'd213: 64'b0001001000111011000011011011011000000010011101111010101001011010;
		8'd214: 64'b1000100100001001001010001110000000100100000000110010000010011000;
		8'd215: 64'b0110101111000111100000101010011001100001111100110101111000101011;
		8'd216: 64'b1111010000101010100101000111001010011010000110001100010001010111;
		8'd217: 64'b0100000100011110111101011101000011010100001001111001010000010100;
		8'd218: 64'b0010001010110110000011100011010000000000000111111101010001000101;
		8'd219: 64'b0101100100011000000000000011100000101001110011011100000001011001;
		8'd220: 64'b1001000001011000001100100011011010000000000011000110100000011001;
		8'd221: 64'b1000000110001101000100000100001010010100000110010001000000000111;
		8'd222: 64'b0110101001111010100011100000101101101010010111101111001001000000;
		8'd223: 64'b0000011010111000100010011000010010000111100100010001100010000000;
		8'd224: 64'b0010011111100001101101101010000000000010011000001011101110100011;
		8'd225: 64'b0010011010000000100100100000110010100001101000100010001010010100;
		8'd226: 64'b0100101101011011101010010000000101001000010100100100010100000010;
		8'd227: 64'b1000111001000110010111001000101000001100100111100100101111101001;
		8'd228: 64'b1001101110001100000000111000101000011001110110000010000111011000;
		8'd229: 64'b0001000010100100000111100000000100100001000011001010111000010000;
		8'd230: 64'b0001001001001011010010010001001010000011000001111000001110001011;
		8'd231: 64'b0101100100101100001010101011010101101000011010100000101010101110;
		8'd232: 64'b0010001000000000100001101111100111001010101001101110010011100100;
		8'd233: 64'b1000110010101001110010001010001010011010011011001000001010100000;
		8'd234: 64'b0011101011000100010101000001000000110011100000010101101011001010;
		8'd235: 64'b0110100101000000111100100011010010001011010001100001100000100000;
		8'd236: 64'b0100100100011000010101100011000011101101101100101100000001011011;
		8'd237: 64'b0100100001100000000000101011011011011110011011110100000110101000;
		8'd238: 64'b0110010011011001101110000100010010001011010000110110001010001001;
		8'd239: 64'b1000100000001000110110110000100010001001100000011001011101100100;
		8'd240: 64'b0101001000100000010000110101001011010001010000110100100100111001;
		8'd241: 64'b0000000001001011110000101010100110000100010111110100000000011110;
		8'd242: 64'b0000000111100111010000000001100000100000001001110001010010011010;
		8'd243: 64'b0001011001100010010000100010001100111011001011101111011000100111;
		8'd244: 64'b1110000100011101011110000101000001000111110001010011011001111000;
		8'd245: 64'b0000100001010000100001000100000010000101101111010000000010010100;
		8'd246: 64'b1000100100000001010101011001001000100100010000001101000100001010;
		8'd247: 64'b1000010100100110001101110011010100001110101101000100001010011001;
		8'd248: 64'b0110111000101010001000000101011100100111000000010110101101011000;
		8'd249: 64'b0111110000110011000001001011000010000101101100000101001000011001;
		8'd250: 64'b0100100000000011000001000100101000110100110010000000110001000010;
		8'd251: 64'b0000010001100111100100000010110101000001110001000100010000000110;
		8'd252: 64'b1001000100000110110110000010100001101001000101001011000000100101;
		8'd253: 64'b1001101100001010100000000101111111000011010111100010011100101101;
		8'd254: 64'b1001110010011001100111001110001111111100101110101001011001000110;
		8'd255: 64'b1000000010001000111010011000000000100010011001001000100011011010;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page3(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1001011001111000101111100110010111000000101101001011010101100011;
		8'd1: 64'b0001011110100111110101100110111101100100101101010110111110111111;
		8'd2: 64'b1111111110010100000011101001001110110101100101100000011110011111;
		8'd3: 64'b1001001000011000111111000011011010010100000100000010010000010010;
		8'd4: 64'b1111000001100100010100010111100011100000110011010010011001111100;
		8'd5: 64'b0011010010100001110001110101010001111101001011011111101111111100;
		8'd6: 64'b1101100101100000100000110001100001101001011010101110101101101000;
		8'd7: 64'b0000011101010001010011000000110000101110000011100010000110000000;
		8'd8: 64'b1011111011011111001100010001000000101001001111100011101100011110;
		8'd9: 64'b1110101010000000000011010000101110001011000010101010011100010101;
		8'd10: 64'b0100001001011010010101100111101000000010011110001110000011111000;
		8'd11: 64'b0110100011011000010000001110101100001100011011100110111101111111;
		8'd12: 64'b0100110011111010100011101010011101001010110111101001101000110111;
		8'd13: 64'b1111100111000010010111001100010010011000000100000101101101000001;
		8'd14: 64'b0001001100110010000110110110011101010010110100100011010000111101;
		8'd15: 64'b1111010010000100001010001010000001110110000111010000110001100011;
		8'd16: 64'b1101100111011100101001011101000111100000100010101010110001010001;
		8'd17: 64'b0001001100101100010010000100000110100001001011011100000010100001;
		8'd18: 64'b0101111010010111001110111100111101010111100101100101101100001000;
		8'd19: 64'b0111100100010011011000111001001110011001011011011101001100011100;
		8'd20: 64'b1010000010111000101110001110101110001101101011001011111000101010;
		8'd21: 64'b1001101011100010101010111110001110100110110000101010111011001101;
		8'd22: 64'b1101100000110010110011001010101011000100110111101000110010001011;
		8'd23: 64'b0110000000111101110010000111111101100001101110011100111101111111;
		8'd24: 64'b1000111000001100100000011000100111101100101111001110111011100111;
		8'd25: 64'b0111001010001001111011111011010001101010000001010001001010000010;
		8'd26: 64'b0101010001000101101000101000010010001010101010000100101111001000;
		8'd27: 64'b1100111101011110110111110101011011001011111101110110100101011100;
		8'd28: 64'b1010101000101100001101111111010101110010101011100010111011001100;
		8'd29: 64'b1001100111010011100011010010011110001111110001001000111001101001;
		8'd30: 64'b0001010110000010010001110101001001100011011001100100001010001000;
		8'd31: 64'b0001100100010110010001011101100001110000000010000100001010101011;
		8'd32: 64'b1111111111101010000110111101100010111111110001111100100001010100;
		8'd33: 64'b1011001001011111101111010100001101101110100101011110100000100101;
		8'd34: 64'b0101110110000111100011111110011001100011100101100001011110100010;
		8'd35: 64'b0000010101000011010100110010000111001111110010010001001100101100;
		8'd36: 64'b1100010000000000101000111101110100011011010011000111001011001101;
		8'd37: 64'b0110100001000100101010011110000010111000101010010011010110110000;
		8'd38: 64'b1111110001111001100001110100001001001111011000011001011100000011;
		8'd39: 64'b0011001010111110100101001000110110110111110111101111001100001001;
		8'd40: 64'b0101111101000011000001101110101101111010100000110010011010010111;
		8'd41: 64'b1001100100010110000010000111101100001010110001101000101100001100;
		8'd42: 64'b1000001011111100011110111000101010111000011010000110011101001001;
		8'd43: 64'b1011110111001100111011100111010010011101001101101011010000100100;
		8'd44: 64'b1100011000000001000010110101001111000010010010001111101010011011;
		8'd45: 64'b0111100101010110110111010000001101110111010011111101100000101010;
		8'd46: 64'b1000000000101001001010011101111110001100001111001000101101001110;
		8'd47: 64'b0111010101010010100000100110000101110101000011000010011000001000;
		8'd48: 64'b1000011111101000101000100100010100101000010111110010100100001101;
		8'd49: 64'b0111100001001001000110111110000100011010010000111000101100110010;
		8'd50: 64'b0001111001011001110111110110110111111110110011011001111011011011;
		8'd51: 64'b1111111110000110101001100111001111100001110000010110110110111000;
		8'd52: 64'b1101110001000001101111100000100101111001011001010100000001011001;
		8'd53: 64'b1011100011000101011111100100001001111000011101110011100111101111;
		8'd54: 64'b0000011110110110111001100111011000100110000101101010011001111100;
		8'd55: 64'b1000110111100110010000011001001110011000100110110000011111110111;
		8'd56: 64'b1100001001001000101011000000001000001010001001010010010010001010;
		8'd57: 64'b0001000011111101010000100100000001011010011010001110000100000011;
		8'd58: 64'b1000000111100100110100001100001010010100010100101101100001100110;
		8'd59: 64'b0010011001011001001001110110000001100110011111010011010100110010;
		8'd60: 64'b1010011000111111011100101111111100011100011011100001101011111111;
		8'd61: 64'b0110101000111000011000000011000111111110111010110010110011010110;
		8'd62: 64'b1100011010101000101101010101100111100010111001011001011101011111;
		8'd63: 64'b1011000010001100110100001001111101101010000100000001100101001001;
		8'd64: 64'b1110011100100011001000110011001110110110111000110001011111110011;
		8'd65: 64'b0011100010010110111000000011100000010110111101001101000011111100;
		8'd66: 64'b1110001011011010101110000101111110110000111011110010000011010101;
		8'd67: 64'b0011111000110001000011111011110010010011010100001000101011011010;
		8'd68: 64'b1010010011100101001001001000001010000100110010111100010110001000;
		8'd69: 64'b1101100000000001100000000011101000001101101010111001100000000010;
		8'd70: 64'b1000110110010000000010101001111010011000010100011000100011111110;
		8'd71: 64'b0010010111001110000000111000111000101100011011000010111010001110;
		8'd72: 64'b0000011111001011101100111001000000101011101001111000001111000110;
		8'd73: 64'b1111101010000000000110001100010101110011111011110001101001000011;
		8'd74: 64'b0011011111110111011011101110011111111110011100001101111110110101;
		8'd75: 64'b0100100101001011000011110001101100101001000110001000100001001001;
		8'd76: 64'b1000100011010100000101001101010001001100111101011001010010110110;
		8'd77: 64'b1101100010010011110000010110111011111100110100111100100111100111;
		8'd78: 64'b1111100111011100110011000101110011101100100011001111110000001101;
		8'd79: 64'b1000011110100001111110100001101100100100000010110111010000010001;
		8'd80: 64'b1111010110110100000101000101011011110111010101100010011100110010;
		8'd81: 64'b1000010111111011010001111010100101000101011010110110110110001101;
		8'd82: 64'b1110000110100000111011011001001000010111100001001001010000010000;
		8'd83: 64'b1000001110001111111011010000110010111100101010101110000100101110;
		8'd84: 64'b0110001111101111111111110011110101100001011101000100101010001100;
		8'd85: 64'b0000111000100111001100000110011000101010111101000010111111100100;
		8'd86: 64'b1010010001001110001111100110010100101101010001011111110101001101;
		8'd87: 64'b1111100010100100110001011010000100101000011011100010000000001010;
		8'd88: 64'b1010001111101010111110010001111010100100111011111110111000001110;
		8'd89: 64'b0100010000110000110100010101010000011100111000011010010101101000;
		8'd90: 64'b1101010110110110000010011001100111011011101110100010101101010100;
		8'd91: 64'b0011110101100001010001000011001010111111100000000001000000000110;
		8'd92: 64'b0011010111100011111000001101000100111001000000011011100010010001;
		8'd93: 64'b1010111010001000101001101010100010101101001000000101001001001011;
		8'd94: 64'b0101101011111010100111111011100001011101111101100001101101000010;
		8'd95: 64'b1111010110000011010001010010110000010110101010000110011000011011;
		8'd96: 64'b1011111101011010100111011001001011111011110111101001011110010010;
		8'd97: 64'b1010111000111111110100100001011111101111001001000001110000000001;
		8'd98: 64'b1110000011101011011100110110110101110101011000110101111101101011;
		8'd99: 64'b1011001001110000111010100110111010010100111101000100001101110010;
		8'd100: 64'b0000101100001000100111101010111010011001100000001101111010001111;
		8'd101: 64'b1010110010011111011111101100010101010000001001111011011010001011;
		8'd102: 64'b0011101000011100001100100001010001101010010111100011111010001000;
		8'd103: 64'b1110010011110100101110100101000110111100110100000100011101010100;
		8'd104: 64'b1101011000000011000111110000000010100000101101100101001111011001;
		8'd105: 64'b1111111100101000011010111110110011100110100110010101100100000100;
		8'd106: 64'b0100101101111001010001100100101001111010111000010100001101011010;
		8'd107: 64'b0101010101010111010010100010110111011100000001000110000101011100;
		8'd108: 64'b1010101011100100011001101010101011010010101111100110010010101010;
		8'd109: 64'b1110010100001100110010011010011100010010001010010110100110000110;
		8'd110: 64'b0001110011101011000100000011111010001010111101101011001001110000;
		8'd111: 64'b1101101011000101100110010110011001110001100100111111100100110011;
		8'd112: 64'b0001001000011101110111100000011111010110001110100111110000000011;
		8'd113: 64'b1001000000011011101100001111001111011100000011110001000001010011;
		8'd114: 64'b1011110010001100100001001001110100101011101011010001110110110001;
		8'd115: 64'b0100000110111101011101011100001001110101001110100011000000100110;
		8'd116: 64'b0110001000101101001010010101010010110111000100110011111000111100;
		8'd117: 64'b0000011111110111001110100111000001000111011011110110111111111101;
		8'd118: 64'b1111111100000011010000011001111000011010101010010010001110101110;
		8'd119: 64'b0100111010010110000111110001001011101110100111111000011110010011;
		8'd120: 64'b1000100010110111011000101101011100101011101101010100111010100011;
		8'd121: 64'b0111111011011100111010100110101011010100111110001110001111100000;
		8'd122: 64'b0110001100100101011101000000111000110110111001010110001011100110;
		8'd123: 64'b0100000111100011110110011110100001100000011010111110000101101110;
		8'd124: 64'b0101100000110010100001011011110101000001111000101000000111011010;
		8'd125: 64'b0111100000011000101111000001010101111000111101100010010000110011;
		8'd126: 64'b1010001100111010000101000000101011000111100010101110100110000111;
		8'd127: 64'b0001010101000111111011110110011100000101001001000000001100101101;
		8'd128: 64'b0001110110110110101111010100001101111000010001001100111000010011;
		8'd129: 64'b1001100110011010110111010111000101111001101000010010001101000000;
		8'd130: 64'b1100010100111100100100000101111110011111111001001101011001011111;
		8'd131: 64'b1101110111010001101111011010100011101011110000111101111010101000;
		8'd132: 64'b0111110111111111101110111011000100010001100000101111011110000111;
		8'd133: 64'b1001111100110100101011101101101111011011000110010100011001000001;
		8'd134: 64'b0000110111001011010001111111000111110011101010101110111101001000;
		8'd135: 64'b0111011001111010000000100111100000101111111100110110111011001000;
		8'd136: 64'b1010000011000101100000111110001001101001111010010010010011000110;
		8'd137: 64'b1101011111010101101001111111011110010000111101010001000110100101;
		8'd138: 64'b0111010101010111111100111001110111101100010011110111000001001100;
		8'd139: 64'b0101110010111001101010101111100010000101001011000110100101100111;
		8'd140: 64'b0000101011001100100011011000000101001010110101100000101011011000;
		8'd141: 64'b0100100110111100000110111000111110010100101100000010111110111101;
		8'd142: 64'b1100111100111111111110000011101111101010001111100010101011110101;
		8'd143: 64'b1110110111100010000100111110011100111000001111110000001001001111;
		8'd144: 64'b1001010101111101100100011111100010111101100111011001011000110100;
		8'd145: 64'b0011100010110101011001010101110100000110001010000100001101111111;
		8'd146: 64'b0110110111110110011000011110110010101011001101100000100111110101;
		8'd147: 64'b0110100000000100100000101011001110100011101000011101100010010010;
		8'd148: 64'b1000011010000111010100010001100001001000101010000001101000000100;
		8'd149: 64'b0010100101110110000000111111011000011001001011100000101001000110;
		8'd150: 64'b1110100010010100111011000011011111101000110101000111111110110001;
		8'd151: 64'b1101000101110011100111000101100010010100000110001011010101000000;
		8'd152: 64'b1010101000100101111010100111111111111110010111111010111011101111;
		8'd153: 64'b1111011110010001101110111001011011011001101100011011111010110001;
		8'd154: 64'b0110010100101010111010011111001101001101010001011110111101001110;
		8'd155: 64'b0100110100100110110101010010100001111000100001010100110000010000;
		8'd156: 64'b0110000101011101101010110001001000011000011001110111111100011010;
		8'd157: 64'b0111010110001000110100001111000011010011110000000101000111101010;
		8'd158: 64'b0100110101001111010001001010001101100101100010001100010001110010;
		8'd159: 64'b1000110101100110101100101111000010100000011011100010010111101110;
		8'd160: 64'b0111110000010110100000011111000100100101111001000100010101001101;
		8'd161: 64'b1000101000110110111001101011101010101101000100101010010010111010;
		8'd162: 64'b0111011011011001011111011101001000100110010010100100100111101011;
		8'd163: 64'b1111011001111011110001001111101001100101111110010001010010101010;
		8'd164: 64'b1000100100011101000110010010111110001001100000010011001110001101;
		8'd165: 64'b0101111001000101100011111001001100101111110011010100111110011011;
		8'd166: 64'b0001010000011111101111011111111001110101101111011011111111110010;
		8'd167: 64'b1010010011100001101000111100011111101100001000111000101101001010;
		8'd168: 64'b0011101000101000110111001000110110111110001010000001100101011101;
		8'd169: 64'b0101011110001011110111111100000110011100100010001100101110000111;
		8'd170: 64'b0000101100001111101110101110101100001010010011100000100101001010;
		8'd171: 64'b0111110111101100001011101010011101001111011011010000110000000001;
		8'd172: 64'b1010111010101111001010111111100000101001110011111010000001010001;
		8'd173: 64'b0001011111000011000000010100101001000101110000101100001110001010;
		8'd174: 64'b1011011101100110110111100110010001111100100011010111111010111000;
		8'd175: 64'b1011011010011011001110111111101010110010011110111111100010101011;
		8'd176: 64'b0111011100011111011111111111101101010101101101000011110110111011;
		8'd177: 64'b0011100010010111101101000111100000111000100001001011100011010101;
		8'd178: 64'b0010101111000010101001000001100010000101000000100011010100000011;
		8'd179: 64'b1110110011100110111111111011011111111111111000101110011001110110;
		8'd180: 64'b1011001000000010101100010000001010011010000111000000010001100011;
		8'd181: 64'b1101000110010010011110001110011011011001001010100110100010010110;
		8'd182: 64'b1100000011111000010010111001101000101011111110100010100110001000;
		8'd183: 64'b0111000010111000001111000000100000011011111111101111010110001100;
		8'd184: 64'b0110100100101111001111101000010101001111000001101011101011000000;
		8'd185: 64'b1001010100011001011010000000101001001100010101000101100111000101;
		8'd186: 64'b1101001101110111010010001101101111011000000101000100000101111011;
		8'd187: 64'b1101010101101011001011010000100011101101001001010001111110001111;
		8'd188: 64'b0010001010001000010111011101100000001100110010100001111001001101;
		8'd189: 64'b0110100010010011100100000100011001100000010100101100000100101110;
		8'd190: 64'b0001010111110010010101110110010111001110001111101111011001100111;
		8'd191: 64'b1100001001111110111011100001000100110011010010101111101100111011;
		8'd192: 64'b1110011101001101111101111110101101000111010010110101010001101000;
		8'd193: 64'b0101010001101101011101111000111001111111000010100011111001000011;
		8'd194: 64'b1101011100110101010100101110000011010111100101010101001101011101;
		8'd195: 64'b1100001000010111110001010001110010000001100100011001110001110100;
		8'd196: 64'b0101000110011001010100010000110001000110110110100101011110111000;
		8'd197: 64'b0011011100100010001101011011100011101110101111100011101100111011;
		8'd198: 64'b0010001000101111110001100010000101100001110011111101010010111101;
		8'd199: 64'b0101111111001111010000000110100101110110110010100101010101100011;
		8'd200: 64'b0101001110010001110110010011100000011100010100101101110010000110;
		8'd201: 64'b1101001001010000111100001011000110010000000100101111011000000010;
		8'd202: 64'b1010100110101110011010110010100000101000111101011110101000110011;
		8'd203: 64'b0110011010101110000001110100111001100111000001100011011111111100;
		8'd204: 64'b1111110010100010100100111000010111101110110110101001001010001100;
		8'd205: 64'b0100011010100100011110110000000110011100011000111010000010011100;
		8'd206: 64'b0101100110000001111111101011010101011000101000010110110110110000;
		8'd207: 64'b0010111000101011101101110110001001101110110010111011011101001010;
		8'd208: 64'b1001101111001001001101110011001111110001010100011011010001000011;
		8'd209: 64'b1001000110111110000010110100010111010000010110100000000100010101;
		8'd210: 64'b1010110000111101111011010101111111100010111111111000100011011010;
		8'd211: 64'b0101011011101101100110101011111111111110010110110101110110111111;
		8'd212: 64'b1000011001000000110101111110111010100110101010110100001101000101;
		8'd213: 64'b0001001000111011001011011011011000010110111111111010101001011111;
		8'd214: 64'b1000100100101101011010011111000100110100000100110110010010011010;
		8'd215: 64'b0110101111000111100000101010011001101011111100111101111011101011;
		8'd216: 64'b1111010000111010100101000111101010011010001110101100010001110111;
		8'd217: 64'b1100100100011110111101011111100011010100001101111011010000011110;
		8'd218: 64'b0111001010110111100111100011010000110010000111111101011001000111;
		8'd219: 64'b0101100100111000010111000011100100101001110011011100000001011011;
		8'd220: 64'b1011000001011000001100100011011010000000010011000111100000011001;
		8'd221: 64'b1000000111001101000110010101001010110101010110010011000001100111;
		8'd222: 64'b1110101101111010101111100000101101101010010111101111001001000011;
		8'd223: 64'b0000011111111010111010111000010010000111100100010011100010000010;
		8'd224: 64'b0011111111101001101101101110000000010010011000011011101111100011;
		8'd225: 64'b0010011010001000100100100000110010100001101000100010001010010100;
		8'd226: 64'b0100111111011011111011010000011101001000010110100101010100000010;
		8'd227: 64'b1010111001010110110111001000111110001100100111100100111111101001;
		8'd228: 64'b1001101110001100000100111000101010011001110110000010000111011000;
		8'd229: 64'b0001010010100100000111101000000100100001000011001110111000010000;
		8'd230: 64'b0001001111011011011010010001011010100011000011111000001110101011;
		8'd231: 64'b0101101100111110101011101011110111111000011010100010111010101111;
		8'd232: 64'b1010011001001110101011101111100111101011111011111111010011101100;
		8'd233: 64'b1010110110101001110010011010001010011010111011001010001010100000;
		8'd234: 64'b1011111011010101011101001001100010110011100000010101101011001010;
		8'd235: 64'b0110100101000001111100100111010010001011010001100001100001100000;
		8'd236: 64'b0100100110011000010111100011000011101101101101101100100001011011;
		8'd237: 64'b0100100001100100010001101011011111011111011011110101010111101000;
		8'd238: 64'b0110010011011001101110000100010110011011010000110110001011101001;
		8'd239: 64'b1000110011101000111110110001100110001001100010011001111101100101;
		8'd240: 64'b0101011100100100010000110101001011110001010100111100100100111001;
		8'd241: 64'b0001000011101011110001101010110110010110110111110100001000011111;
		8'd242: 64'b0000000111111111010000000001100000100000001011110001010011111010;
		8'd243: 64'b0101011001100010110000100010001100111011001011101111011000100111;
		8'd244: 64'b1110000100011101111110001111010101100111111001010011011111111000;
		8'd245: 64'b0010100101011000100001000100100010000101111111010000010010011110;
		8'd246: 64'b1000100100000011011101011011001000100100010100001101000101011011;
		8'd247: 64'b1011010110100110001101110011010110011111111111010110101011011001;
		8'd248: 64'b0110111000101010011010000101011110100111000000010110101101011100;
		8'd249: 64'b1111110100110011000011001011101010000101101100100101001100011001;
		8'd250: 64'b0100100000000011000111100100101000110101111010010001110001001010;
		8'd251: 64'b0100010011100111100100000110110111100101110001000101011000100110;
		8'd252: 64'b1001100110100110110110000010100011101001000101101011001000101101;
		8'd253: 64'b1101101101101110100101000111111111000011011111100011111110101111;
		8'd254: 64'b1001110010111001110111101110001111111100111111101001111001001110;
		8'd255: 64'b1001000010101000111110011100101110100010011001001000100111011010;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page4(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1001011101111000101111100111010111000100101101001011010101110011;
		8'd1: 64'b1001011111100111110111101110111111110110111101110110111110111111;
		8'd2: 64'b1111111110010110000011101001001110110101100101100010011110011111;
		8'd3: 64'b1001101000011000111111001011011010010100000100000010010000010010;
		8'd4: 64'b1111000001100110010100010111100011110000111011010110011101111100;
		8'd5: 64'b0111010011110101111001111101010001111101101011011111111111111100;
		8'd6: 64'b1101100101100010100000110001100001101001011010101110101101101000;
		8'd7: 64'b0000011101010001010011000000110000101110000011100010000110000000;
		8'd8: 64'b1011111111111111101100010001000000101001001111100011101100011111;
		8'd9: 64'b1110101010000010000011010000101110001011100010101010011100010101;
		8'd10: 64'b0100001001011010010101100111101011000010011110001110110011111000;
		8'd11: 64'b1111100011011000010010001110101100001101011011100110111101111111;
		8'd12: 64'b0100111011111010100011101011011101001010110111101001101000111111;
		8'd13: 64'b1111101111000010010111001100010010011110000100000101101101000001;
		8'd14: 64'b0001001100110010000111110110011101010011110101100011010100111111;
		8'd15: 64'b1111010010000100101011001010000001110110000111010101110001101011;
		8'd16: 64'b1111100111111100101001011101000111100011100010101010110001010011;
		8'd17: 64'b0101001100101100010010101100000110101001011011111100000010100001;
		8'd18: 64'b1101111110010111001110111110111101010111100101101111101100001000;
		8'd19: 64'b0111100100010011111101111011001111011001011011011101001100011111;
		8'd20: 64'b1010100010111000101111101110101111001101101011001011111010101010;
		8'd21: 64'b1001101011100010101010111110001110100111110000101010111011101101;
		8'd22: 64'b1101100001110110110011001010101111000100111111101100110010101011;
		8'd23: 64'b0110000010111101110011100111111101100011101110111110111101111111;
		8'd24: 64'b1001111000001100110011011000100111101100101111001110111011100111;
		8'd25: 64'b0111101110001001111011111011010101101010000001010001001010000010;
		8'd26: 64'b0111010001000101111000101100010010001010111011000100101111001100;
		8'd27: 64'b1100111101011110111111110101011011001011111101110110100101011100;
		8'd28: 64'b1110101000101110001111111111110101111110101011110010111011111110;
		8'd29: 64'b1011100111010111100011010010011110011111110001001001111001101001;
		8'd30: 64'b0101010110010010010001110101001001101011011001100100001111001000;
		8'd31: 64'b0001100100010110110001011101100011110001000010010100001010101011;
		8'd32: 64'b1111111111101010000110111101100010111111111001111110101011011100;
		8'd33: 64'b1111001001011111111111010100011111101110100101011110110000100101;
		8'd34: 64'b0111111110000111100011111110011011100111100101110101011111100110;
		8'd35: 64'b0000110101000011010100110010000111001111110110010001001100111100;
		8'd36: 64'b1100010001000100101000111101111100011011010011011111001011001101;
		8'd37: 64'b0110100001000100101110011111001010111000101011010011010111110000;
		8'd38: 64'b1111111101111001100001110100001001001111011100011001011101000011;
		8'd39: 64'b1011001011111110110101011010110110110111111111111111011100001101;
		8'd40: 64'b0101111111000011000001101110101101111010100000110010011011111111;
		8'd41: 64'b1001101100010110000010100111101100001010110001101000101100001100;
		8'd42: 64'b1000101011111100011110111010101010111000011010100110011101001001;
		8'd43: 64'b1011110111001100111111100111010110011101001111101011010000110100;
		8'd44: 64'b1100011000010001000010110101001111000010011010001111111011011011;
		8'd45: 64'b0111101101010110110111010000001101110111010011111101110000111011;
		8'd46: 64'b1000100000101001001010011101111110001100001111001000101101001111;
		8'd47: 64'b0111010101110010101000101111000101110101000111000010011000001000;
		8'd48: 64'b1100011111101001101000110100010100101011010111111111100101001101;
		8'd49: 64'b1111100101001001010110111111000100011010010000111001111110111110;
		8'd50: 64'b0001111001011001110111111110110111111110110011011001111011011011;
		8'd51: 64'b1111111110000110101001100111101111110011110000010110111110111000;
		8'd52: 64'b1101110001000001101111110000100101111011111001010100000001011001;
		8'd53: 64'b1111100011000101011111100101011111111001011101111011110111101111;
		8'd54: 64'b0000111110110110111001100111111000100110000101101010111001111100;
		8'd55: 64'b1000110111101110010000111001101110011000100110110100011111110111;
		8'd56: 64'b1100001001001000101011000000001000001010011001010010010010001010;
		8'd57: 64'b0001100011111101010000100101000101011010011010011110000100000011;
		8'd58: 64'b1100000111100100110110001100101010010100010101101101100101100110;
		8'd59: 64'b0010011001011001001001110110000001100110011111010011111100110010;
		8'd60: 64'b1011011000111111011101111111111110011100011011100011101011111111;
		8'd61: 64'b0110101000111101111001001011000111111111111010110010110111011110;
		8'd62: 64'b1100011011101000101101010101101111100010111011011001011101011111;
		8'd63: 64'b1011100010001100110110001011111101101110100110100001111101001001;
		8'd64: 64'b1111111101101011001001110011001110110111111100110011011111110011;
		8'd65: 64'b0011100010010111111000000011100010110110111101001111000011111110;
		8'd66: 64'b1110101011011010101110000101111111110000111011110010000011010101;
		8'd67: 64'b0011111000110001000011111011110010110011110100001000101011111010;
		8'd68: 64'b1010010011100101001001001000101010000100110010111110010110001000;
		8'd69: 64'b1101100000000001100000000111101000001111101010111001100000000010;
		8'd70: 64'b1001110110010100000010101111111010011000010100011000100011111110;
		8'd71: 64'b0010110111001110000000111000111000101100011011000010111010001110;
		8'd72: 64'b0100011111001011111110111001100000101011101001111000001111100110;
		8'd73: 64'b1111101010000100000111001110010101110111111011110001101001100111;
		8'd74: 64'b0111111111110111011011101110011111111110011100001101111111111101;
		8'd75: 64'b1101100101001011010011110001101100101001000110101000111101001001;
		8'd76: 64'b1101100011010110010111101101110011001100111101011001010011110110;
		8'd77: 64'b1101100010010011110000111111111011111101110100111100100111100111;
		8'd78: 64'b1111110111011100110011101101110011101100110011001111110000011101;
		8'd79: 64'b1010011110100001111110100001101100100101000010110111010000010001;
		8'd80: 64'b1111011110110100101111000101011011110111010101100011011100110010;
		8'd81: 64'b1100011111111011010001111010100101001111111010110110110110101101;
		8'd82: 64'b1110000110100100111011011101001000010111100001001001010010010000;
		8'd83: 64'b1010001110001111111011110000110010111100111010111110100110101110;
		8'd84: 64'b0110011111101111111111110011110101100001011101000100101110011100;
		8'd85: 64'b0010111101100111001100100110011001101010111111110010111111100100;
		8'd86: 64'b1110110001001110001111100110011100111101010001011111111111101101;
		8'd87: 64'b1111100010101100110001011110010100101110011011101010000010001011;
		8'd88: 64'b1010001111101010111110010001111010100110111011111110111100011110;
		8'd89: 64'b1100010000110000110100110101110000011100111000011110011101101100;
		8'd90: 64'b1101010110110111000010011001100111011011101110101010101111010100;
		8'd91: 64'b0011110101100001011001000011001010111111110000000101000000100110;
		8'd92: 64'b0111010111100111111000001101000100111001010000011011100010010001;
		8'd93: 64'b1010111010001000101011101010100010101101101010000101001001001011;
		8'd94: 64'b0101101111111011100111111011100001011101111101100001101101000010;
		8'd95: 64'b1111010110000111010001010010110000010110101010010110011000011011;
		8'd96: 64'b1011111101011010100111011001001011111011110111101001011110010011;
		8'd97: 64'b1010111100111111110110100101011111101111001001000001111000000001;
		8'd98: 64'b1110000111111011011100110110111101110111011010111101111101101011;
		8'd99: 64'b1011001001110000111010100111111010010111111101000110001101110010;
		8'd100: 64'b0000101111001000100111101010111010011001100010001111111010101111;
		8'd101: 64'b1110110010011111111111101100010101010000101011111011011010001111;
		8'd102: 64'b0011101010011100001110100001010001111110010111100011111010001000;
		8'd103: 64'b1110010011110110101110100101000111111110110100000100011101010100;
		8'd104: 64'b1111011000000011000111110001000110110011101101110101001111011011;
		8'd105: 64'b1111111110101000011010111110110011100111100111010101110100000100;
		8'd106: 64'b0100101101111011010001100100101001111010111000010100001101011010;
		8'd107: 64'b0101010101010111010010100010111111011100100011000110001101011110;
		8'd108: 64'b1010101011101100011001101010101011110010101111100110010010101010;
		8'd109: 64'b1110010100001100110010011010011100010010001010010110100111000110;
		8'd110: 64'b0101110011101011000100000011111010001010111101101011001001110000;
		8'd111: 64'b1101101011000101110110010110011001110001100100111111100100110011;
		8'd112: 64'b0001011000011101110111110010011111011111001110110111110000100011;
		8'd113: 64'b1001000000011011101100001111001111011100000111111001000001010011;
		8'd114: 64'b1011110010001100100011001001110100101011101011010001110110110001;
		8'd115: 64'b0100000110111111011101011100101001110101011110100111000000100110;
		8'd116: 64'b0110011000101101001010010101011010110111000100110111111000111110;
		8'd117: 64'b0011011111110111001110100111001001100111111011110110111111111101;
		8'd118: 64'b1111111101001011010000011001111011011010111010010010001110101111;
		8'd119: 64'b0100111010110110100111111001001011111110100111111000111110010111;
		8'd120: 64'b1000100110110111011010101101011100101011111101110100111010100011;
		8'd121: 64'b0111111011011100111010100110101011010100111110001110001111100000;
		8'd122: 64'b0110111100100101011101000010111001110110111001110110001011100110;
		8'd123: 64'b0110000111100011110110011110110011100000011110111110000101101110;
		8'd124: 64'b0101100000110010100001011011110101010001111000101000000111111110;
		8'd125: 64'b0111101101011000101111000001010101111000111101100010010101110011;
		8'd126: 64'b1010001100111110100111000010101011000111110011101110101110000111;
		8'd127: 64'b0001010101100111111011110110011100000111001001000010011100101101;
		8'd128: 64'b1001110110110110101111010100001111111000010111001101111001011011;
		8'd129: 64'b1001110110011011110111011111000101111001101001010010001101100000;
		8'd130: 64'b1100010111111101110100000101111110011111111001011101011001011111;
		8'd131: 64'b1101110111010001111111011010100011101011111000111101111010101000;
		8'd132: 64'b0111110111111111101110111011110100110101100000101111111110000111;
		8'd133: 64'b1001111100110100101011101101101111011011011111011100011001000001;
		8'd134: 64'b0100110111001011010011111111000111110011111010101110111111001000;
		8'd135: 64'b0111011101111011000001100111100000111111111100110110111011011000;
		8'd136: 64'b1110010011000101100001111110001011101011111010011010110011001110;
		8'd137: 64'b1101011111110101101001111111011110010001111101011001000111100101;
		8'd138: 64'b0111010111010111111100111101110111101101010011110111000001001100;
		8'd139: 64'b0101110010111001111010101111100010000101001011001110100101110111;
		8'd140: 64'b0000101011001100110011011000000101001010110101100000101011011000;
		8'd141: 64'b0100100110111100000110111000111110010100101101000010111110111101;
		8'd142: 64'b1110111100111111111110000111111111101110001111110010111011111101;
		8'd143: 64'b1110111111100010000100111110011100111000001111110100001001001111;
		8'd144: 64'b1001010101111101101100011111100010111101101111011001111000111100;
		8'd145: 64'b0011101110111101011001010101110100110110001010100100001101111111;
		8'd146: 64'b1110110111110110011000011110110010101011011101101000100111111101;
		8'd147: 64'b0110110000000100110100101011101110100011101000111101100010010010;
		8'd148: 64'b1000011010000111010100010001100001001000101010000001101000100100;
		8'd149: 64'b0011101101110110100010111111011110111001011111100000101001100110;
		8'd150: 64'b1111100010010110111011010011011111101000110101010111111110110111;
		8'd151: 64'b1101010101110011100111000101100010010110001110001011010111000100;
		8'd152: 64'b1110101000100111111010100111111111111110010111111010111111101111;
		8'd153: 64'b1111111110010001101110111001011111111011101110011111111010110001;
		8'd154: 64'b0110010101101010111011011111001101001101010011011110111101001110;
		8'd155: 64'b1100111100110110110101010010100001111100100001110101110000010100;
		8'd156: 64'b0110000101011111111010110001001000011001011011110111111100111010;
		8'd157: 64'b0111010110001000110100001111000011010011110000001101000111111010;
		8'd158: 64'b0110110101011111011001101110001101100101100011001100010001110010;
		8'd159: 64'b1001110101100110101100101111001010100000011011110010010111111110;
		8'd160: 64'b0111110100010110100000011111010101100101111011010100010101001101;
		8'd161: 64'b1010101000110110111001101011101010111101000101101110010110111010;
		8'd162: 64'b1111111011011011011111011101101000100110110010100100100111101011;
		8'd163: 64'b1111011001111011110101001111101001100101111110111001010010111010;
		8'd164: 64'b1001100100011101000110010011111110001011100100111111001110001101;
		8'd165: 64'b0101111011000101100011111001101100101111110011011100111110011011;
		8'd166: 64'b0001010100011111111111011111111011110101101111011011111111110011;
		8'd167: 64'b1110010111100011101000111100011111101101101000111000101111001010;
		8'd168: 64'b0011111000101000110111001100110110111110001010111001110111011101;
		8'd169: 64'b1101111110001111110111111100010111011100100010011100101110011111;
		8'd170: 64'b0100111100001111101110101110101100001010110011100000100101001010;
		8'd171: 64'b0111110111101100001011101010011101011111011011010000110000000001;
		8'd172: 64'b1110111110111111001010111111100001101011110111111010110001110001;
		8'd173: 64'b0011011111000011000000111100101001001101111000101100001110001010;
		8'd174: 64'b1011111111100111110111100110110001111100100111010111111010111001;
		8'd175: 64'b1011011011111011101110111111101010110010111110111111100011101011;
		8'd176: 64'b0111011100011111011111111111101101110101101111010111111110111011;
		8'd177: 64'b0011101011010111101101000111100000111000100001001011100111110101;
		8'd178: 64'b0010101111100010101001100001100010110101000000100011010100000011;
		8'd179: 64'b1110110011100110111111111011011111111111111001101110011001110110;
		8'd180: 64'b1011001100100010101100010000011110111010010111001100010001100011;
		8'd181: 64'b1101000110110010011110001110011011011001001010100110100011110110;
		8'd182: 64'b1100100011111000010010111001111000101011111110100010100110001000;
		8'd183: 64'b0111010010111000001111000010100100111011111111111111011111001100;
		8'd184: 64'b0110100100101111001111101000010101001111000001101111101111010000;
		8'd185: 64'b1001010101011101011010000010101001011100010101101101100111000101;
		8'd186: 64'b1101001101110111111010001101101111011000010101000100000101111011;
		8'd187: 64'b1101010101101011001011010001100011111101001001010001111110001111;
		8'd188: 64'b0111001010001010010111011101110010011100110011100001111001001101;
		8'd189: 64'b0110101010010011101100010110011001100000010100101100010110101110;
		8'd190: 64'b0001010111110010010101110110010111011110001111101111011001100111;
		8'd191: 64'b1100101001111110111011100001000100111011010010101111101100111011;
		8'd192: 64'b1110011101001111111101111110101111100111011011110101011001101000;
		8'd193: 64'b0111010001101101011101111000111001111111000010110011111101000111;
		8'd194: 64'b1101011100110101010100101110000011010111110101011101001101011101;
		8'd195: 64'b1100101000010111110111010001110010000001100100011001110001111101;
		8'd196: 64'b0111000110011001010100010000110001000110110110100101011110111000;
		8'd197: 64'b0011011100100010001101111011101011101110101111100011101100111011;
		8'd198: 64'b0010101000101111110001110010110101100011110011111101010011111101;
		8'd199: 64'b0111111111001111011000001110101111110110110011100101010101100011;
		8'd200: 64'b0101011110010001110111010011100000011100110100101101110010110110;
		8'd201: 64'b1101001001010010111100001011000110010001000100111111011000100010;
		8'd202: 64'b1010100110101110011010110010100000101000111101011110101000110011;
		8'd203: 64'b0110011010101110100101110100111001100111100001100011011111111111;
		8'd204: 64'b1111110010100010100100111010010111101110110111101001001010001110;
		8'd205: 64'b0100011010110101011110110000000110011100011000111011000010011100;
		8'd206: 64'b0101100110000001111111101011010101111000101010010110110110110000;
		8'd207: 64'b0010111111101011101101110110001001101110110010111011011101001010;
		8'd208: 64'b1001101111001011101101110011001111111011010110111011010001000011;
		8'd209: 64'b1101000110111110100010110101010111010001010111100000010101010101;
		8'd210: 64'b1111110100111101111011010101111111101010111111111000100011111111;
		8'd211: 64'b1111011011111111100110101011111111111110010111110101110110111111;
		8'd212: 64'b1000011101000010110101111110111010100110101010110100001101000101;
		8'd213: 64'b0001111000111011001011111011011000010110111111111010101001111111;
		8'd214: 64'b1000100100111111011010011111000100110100000100110110010010111010;
		8'd215: 64'b1110111111000111101100111011011101101111111100111101111011101011;
		8'd216: 64'b1111010001111010100111000111101010011010001111101101010001111111;
		8'd217: 64'b1101100100011110111101011111110011010100001111111111010000011110;
		8'd218: 64'b0111001010110111100111100111011001111010000111111111011001000111;
		8'd219: 64'b0111100100111001010111000111100100101001110011011100110001011011;
		8'd220: 64'b1011000001011100001100100011111010000000010111000111100010011001;
		8'd221: 64'b1011000111101101001110011101101010110111010110010011000001100111;
		8'd222: 64'b1110101101111010101111101000101101101010010111111111001011000011;
		8'd223: 64'b0001111111111010111110111000010010000111100100011011100010000110;
		8'd224: 64'b0011111111101001101101101110100010010110011010011011111111101011;
		8'd225: 64'b0110011010011100100110100000110010100001101000100010111010010101;
		8'd226: 64'b1110111111011011111011010001011101001100011110111101010101001110;
		8'd227: 64'b1110111001010110110111001100111111001100110111100100111111101101;
		8'd228: 64'b1011101110011100000110111000111010011001110110000010000111011001;
		8'd229: 64'b0011010010100100001111101000000100100001010011001110111001010000;
		8'd230: 64'b0001001111011011011010010001011110110011000111111000001110101011;
		8'd231: 64'b1101101100111110101011111011110111111000011010100010111010101111;
		8'd232: 64'b1011011001101110111011101111110111111111111011111111011011101100;
		8'd233: 64'b1010110110101001110010011010001010011010111011001010001110101000;
		8'd234: 64'b1011111011010101011101001101100010110011100000010101111011011010;
		8'd235: 64'b0111110101000001111100100111010010011011010001100001100001100000;
		8'd236: 64'b0100100110011001010111110011000011101101101101101100110101111011;
		8'd237: 64'b0100110101101100010001101011011111011111011011110101010111101000;
		8'd238: 64'b0110010011011101101110000101011110111011110000110110001011101001;
		8'd239: 64'b1010110011111100111110110101110110001001100010011001111101110101;
		8'd240: 64'b0101011101110100010100110101001011111001010100111100100100111001;
		8'd241: 64'b0101000011111011110011101010110111010111110111110101001010011111;
		8'd242: 64'b0000000111111111010000000001100000100000001011110001010011111010;
		8'd243: 64'b0101011011101011110001100010001100111011001011101111011000100111;
		8'd244: 64'b1110001101011101111110001111010101100111111011011011011111111010;
		8'd245: 64'b1010100111111000100001000100100011000101111111010000010010011110;
		8'd246: 64'b1100110101000011011101011011101010110100010101011101000101011111;
		8'd247: 64'b1011111110100110101101110011010110011111111111010110101011011001;
		8'd248: 64'b0110111000101010111010000111011111100111000000110110101101111100;
		8'd249: 64'b1111110100110011000011001111101010000101101100100101001100011011;
		8'd250: 64'b0100100000001011000111100100101000110101111010010001110011001010;
		8'd251: 64'b1100011011100111110100000110110111100101110001000101011000110110;
		8'd252: 64'b1101100111100110111110000010100111101101000101101111101001101101;
		8'd253: 64'b1101101101101111100101000111111111000011011111110011111110101111;
		8'd254: 64'b1001110010111101111111101110101111111101111111101101111001001110;
		8'd255: 64'b1001000011101010111110011100101110100011111101001000110111011010;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page5(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1001011101111001101111100111010111010100111101001011010101110011;
		8'd1: 64'b1101011111100111111111101111111111110110111101110110111110111111;
		8'd2: 64'b1111111110010110001011111101001110110111100101100010111110111111;
		8'd3: 64'b1001111000011000111111001011011010011100000100000010010100010011;
		8'd4: 64'b1111000001110110010100011111101011110000111011010110011101111100;
		8'd5: 64'b0111111011111101111001111111010111111101111011011111111111111101;
		8'd6: 64'b1111101101101011110010110001100001101001011110101110101101101000;
		8'd7: 64'b0000011101010001010011000000110010101111001011100010000110000000;
		8'd8: 64'b1011111111111111101100010001000100101001001111100011101100011111;
		8'd9: 64'b1110101110011010001011110000101110101011100011101010111100010111;
		8'd10: 64'b0110001101111011110101100111101011000110111110101111110011111010;
		8'd11: 64'b1111100111011100010010001110101101001101011011110111111111111111;
		8'd12: 64'b0100111011111010100111101011011101011110110111101101111011111111;
		8'd13: 64'b1111101111000011010111001100010010011110000100001101101101000001;
		8'd14: 64'b0001011100110110000111110110011111010011110101100011010100111111;
		8'd15: 64'b1111010010000101111011001010010001110110100111011111110101111011;
		8'd16: 64'b1111100111111100101001011101110111101011110011101010111001010011;
		8'd17: 64'b0101001100101101010010101100100110101101111011111100001010100001;
		8'd18: 64'b1101111110010111011110111110111101010111100101101111111100001110;
		8'd19: 64'b0111100100010011111101111011001111011001011011111101011101111111;
		8'd20: 64'b1010100010111000111111101110101111001101101011001011111010101010;
		8'd21: 64'b1001101011100010101011111110001110111111110000111010111011111101;
		8'd22: 64'b1111101011110111110011001010101111000100111111101111110110111011;
		8'd23: 64'b0110001010111101110111100111111101101111101110111110111101111111;
		8'd24: 64'b1101111000001110111111011000100111101100111111001111111011100111;
		8'd25: 64'b0111101110101001111011111011011111101010000001010001101010100010;
		8'd26: 64'b0111010001001101111100111100010011001010111011001100101111101101;
		8'd27: 64'b1100111111011110111111111101011011001011111101110110101111011100;
		8'd28: 64'b1110101010101110101111111111110101111110101011110010111011111110;
		8'd29: 64'b1011100111010111100011110010011110011111110001001011111001101001;
		8'd30: 64'b0101111110010010010001110101001001101011011001100101001111001000;
		8'd31: 64'b0111100100010110110101011101100111110001000010011100111010101011;
		8'd32: 64'b1111111111101011000110111101100011111111111001111110101011011101;
		8'd33: 64'b1111101011011111111111010100011111101110100101011110110000100101;
		8'd34: 64'b0111111110101111100011111110011011110111100101110111011111100110;
		8'd35: 64'b0100110101000011010100111010101111001111110111010001001100111100;
		8'd36: 64'b1100010001000101101000111111111100011011010011111111101111001101;
		8'd37: 64'b0110101001100100101110011111001011111000101011010011111111110000;
		8'd38: 64'b1111111101111001100001110100001001001111111100011101011111000011;
		8'd39: 64'b1011001011111110110101011011110111110111111111111111011100001101;
		8'd40: 64'b0101111111000111000001101111101111111110110000111010011011111111;
		8'd41: 64'b1101101100010110000110100111101100001010110001101000101100011100;
		8'd42: 64'b1100101111111100011110111110101010111000011110100110011101101001;
		8'd43: 64'b1011111111001100111111110111010110011111001111111011011010110100;
		8'd44: 64'b1100011001010101000110111101101111001010011010001111111011011011;
		8'd45: 64'b0111101101010110110111010001101101110111010011111101110000111011;
		8'd46: 64'b1000110000111001001010011101111110001100001111001001111101001111;
		8'd47: 64'b0111011101110010101000101111001101110101010111000010011000001000;
		8'd48: 64'b1110011111101001101000110110010100101111010111111111100101011101;
		8'd49: 64'b1111100101111001010110111111000100111010011110111001111110111111;
		8'd50: 64'b0001111011011001110111111110111111111110110011011111111011111111;
		8'd51: 64'b1111111110000110101001100111111111110011111000110110111110111000;
		8'd52: 64'b1101110001011001111111110100100101111011111001010101100001011011;
		8'd53: 64'b1111100011110101011111110101011111111001011101111011110111111111;
		8'd54: 64'b1000111110110110111001100111111000100110000111101010111011111100;
		8'd55: 64'b1000111111101110110100111111101110011000101110110101011111110111;
		8'd56: 64'b1100011001001100101011001000011010001010011011011110010011001010;
		8'd57: 64'b1101100111111101011000111101000101011010011010011110010101000111;
		8'd58: 64'b1101000111100101110110001110101011010101010101101101100101111110;
		8'd59: 64'b0010111001111001101001110110001001100110011111010011111101110010;
		8'd60: 64'b1111011000111111111101111111111110011100011011100111111011111111;
		8'd61: 64'b0110101010111101111011001011000111111111111010110010110111011111;
		8'd62: 64'b1110111011101000111111011101101111100010111011011011011101011111;
		8'd63: 64'b1011100010001101110110001011111101111110101110100001111101001011;
		8'd64: 64'b1111111101111011001001110011001110111111111100110011011111110011;
		8'd65: 64'b0011100010010111111100000011100010111110111101001111000011111110;
		8'd66: 64'b1111101011011111101111000101111111111000111111110010000111011101;
		8'd67: 64'b0011111000110001000011111011110010110011111100001010111111111111;
		8'd68: 64'b1010010011100101001001001000111010000100110010111110010110001000;
		8'd69: 64'b1101101101001001100100000111101000011111101010111001100000001010;
		8'd70: 64'b1001110110110100000010101111111010011000010111111000100011111110;
		8'd71: 64'b0010110111001110000000111000111000101110011011000010111010011110;
		8'd72: 64'b1110011111011011111110111101101000101011111001111000101111100110;
		8'd73: 64'b1111101010000100001111001110010101111111111011110101101001100111;
		8'd74: 64'b0111111111110111011011111110011111111111011100101101111111111101;
		8'd75: 64'b1101100101001011010011110001101100101001000110101000111101001111;
		8'd76: 64'b1101100011010110111111101101111111011100111101011001110011110110;
		8'd77: 64'b1111111010010011110001111111111111111101110100111100100111100111;
		8'd78: 64'b1111110111011100110011101101110011101100110011001111110001011101;
		8'd79: 64'b1010011110101001111111110001101100100101001111111111010000010001;
		8'd80: 64'b1111011111110101101111100111011011110111011101100111011100110110;
		8'd81: 64'b1100011111111011010001111010100101001111111010110110111110101101;
		8'd82: 64'b1110100111100100111111011101011000010111100001101101110111010000;
		8'd83: 64'b1110101110101111111011110000110010111100111010111110111110101110;
		8'd84: 64'b0110111111101111111111110011111101100001011101000100101110011100;
		8'd85: 64'b0010111101100111001100100110011001101110111111110010111111100110;
		8'd86: 64'b1110111101001110001111100110111100111111010001011111111111101111;
		8'd87: 64'b1111100011101110111001011110110100101110011011101010000010001011;
		8'd88: 64'b1010001111101110111110110011111010100110111111111111111110011110;
		8'd89: 64'b1101110010110000110100110101110000011100111100011110011101101100;
		8'd90: 64'b1101010110110111000011111101100111011011101110101110111111010100;
		8'd91: 64'b0011110101100001111001000011101010111111110000000101110000110110;
		8'd92: 64'b0111110111100111111000001101000101111101010000011011100011011001;
		8'd93: 64'b1010111010101000101011101010100010101101111010001101001101001011;
		8'd94: 64'b1101101111111111110111111111101001011101111111100001101101000110;
		8'd95: 64'b1111010110001111010001010111111001010110101011010111111000011011;
		8'd96: 64'b1011111101111010100111111001001011111011110111101001111111110011;
		8'd97: 64'b1010111111111111110111110101011111101111001001000001111100100101;
		8'd98: 64'b1110010111111011011101110111111101110111011110111101111101101011;
		8'd99: 64'b1011111001110000111010100111111010010111111101000110001101110010;
		8'd100: 64'b1001101111001100100111101010111010011001101010001111111010101111;
		8'd101: 64'b1110110010111111111111101110011111010010101011111011011010001111;
		8'd102: 64'b0011101010011101011110100011010011111110110111100011111110001000;
		8'd103: 64'b1111010111110110101110100101001111111110110101000100111101110110;
		8'd104: 64'b1111011000000111000111110001001110110011101101111111101111011011;
		8'd105: 64'b1111111110101100011110111110110011100111110111010101110110000100;
		8'd106: 64'b0100101101111011010001100100101001111011111101010100001101011110;
		8'd107: 64'b1101010101010111010010100010111111011100100111000110001101011110;
		8'd108: 64'b1010101011101100011001101010101011110110101111101110011110111010;
		8'd109: 64'b1110010100001101110010011010011110010011001010010111100111100110;
		8'd110: 64'b0101110011101111000100101011111011011011111101101011011001110000;
		8'd111: 64'b1101101111011111110110010110011001110101100100111111100100110111;
		8'd112: 64'b1001011100011101110111110010011111011111001110110111111001101011;
		8'd113: 64'b1001100000011011101100001111001111011100000111111011000001010011;
		8'd114: 64'b1011110010001101100011001001110111101011111111010001110110111001;
		8'd115: 64'b0100000110111111011111011100101001110101011110100111000000101110;
		8'd116: 64'b0110011100101111001010011101011110110111001100111111111001111110;
		8'd117: 64'b0111011111110111001110100111001001100111111011110110111111111111;
		8'd118: 64'b1111111101001011110000011001111011011010111110110110001111101111;
		8'd119: 64'b1100111010110110100111111001001011111110110111111001111110010111;
		8'd120: 64'b1100101110110111011010101101111100111011111101110110111110100011;
		8'd121: 64'b0111111111111100111010100111101011110100111110001110001111100000;
		8'd122: 64'b0110111100100111011101100010111101110110111001110110101111100110;
		8'd123: 64'b0110000111100111111110011111110011100000011110111110000101101110;
		8'd124: 64'b0101100000110011100001011011111101010001111000101010000111111110;
		8'd125: 64'b0111101101011010101111110001010111111000111101110010010101110011;
		8'd126: 64'b1011001100111110100111101110101011000111111011101110101110000111;
		8'd127: 64'b1011011101101111111011110110011100000111011001010010011100101101;
		8'd128: 64'b1001110110111110101111011100001111111000110111101101111001011011;
		8'd129: 64'b1001110111011011110111011111000101111001101101010010001111100000;
		8'd130: 64'b1101010111111101110100000101111110011111111111011101011101011111;
		8'd131: 64'b1101110111010001111111011010100011101011111000111111111011101000;
		8'd132: 64'b0111111111111111101110111011111101110101100000111111111110001111;
		8'd133: 64'b1001111110110101101011111101101111011011011111011111111001010011;
		8'd134: 64'b0100110111001011010011111111000111111111111010101110111111001000;
		8'd135: 64'b0111011101111011000001100111101000111111111100110110111111111010;
		8'd136: 64'b1110011011001101100001111110101011101111111011011010111111001110;
		8'd137: 64'b1101011111110101101001111111011110010001111111111001000111110101;
		8'd138: 64'b0111010111010111111100111101111111111111010111110111010001101100;
		8'd139: 64'b0101110010111001111011101111100110000101001111101110100101110111;
		8'd140: 64'b0000101011001100110011011000010101001010110101100000111011011000;
		8'd141: 64'b0100100110111100000110111010111110010110101101000010111110111101;
		8'd142: 64'b1110111100111111111111000111111111101110101111111010111011111101;
		8'd143: 64'b1110111111101011000100111110011100111001001111110101001101101111;
		8'd144: 64'b1011010111111101101100011111100010111101101111111001111010111100;
		8'd145: 64'b0111101110111101011001011101111110110110011011100100011101111111;
		8'd146: 64'b1110110111110110111010011110110010101111111111101000110111111101;
		8'd147: 64'b0110111001000101110110111011101110110011101000111101110010010010;
		8'd148: 64'b1100011110000111110100011001110011001000101010100001101000100100;
		8'd149: 64'b1011101101110110100011111111011110111011011111100000101001100110;
		8'd150: 64'b1111100010110110111111011011011111101001110101110111111111110111;
		8'd151: 64'b1101010101110011101111000101101010110110001110011011010111000100;
		8'd152: 64'b1111111011101111111010111111111111111110010111111110111111111111;
		8'd153: 64'b1111111110010011101110111001111111111011101110011111111010110001;
		8'd154: 64'b0110010101101011111011111111001101001111111011111110111101001110;
		8'd155: 64'b1100111100110110110101010010110011111100110001110101110000110110;
		8'd156: 64'b0111001111111111111010110101001111011001011111110111111100111010;
		8'd157: 64'b0111010110011000110100011111010011010011110010001101000111111010;
		8'd158: 64'b0110110111011111011101101110011101101101100011011100010001110011;
		8'd159: 64'b1011110111110110101100101111101010110000011011110011011111111110;
		8'd160: 64'b0111110100010111101001011111110101110111111011010100011101001101;
		8'd161: 64'b1010101000110110111101111011101010111101001101101110010110111010;
		8'd162: 64'b1111111011011011111111011101101001100110110110100100100111111011;
		8'd163: 64'b1111011111111011110101101111101011111101111110111101011011111010;
		8'd164: 64'b1001100100011101000111010011111110001011100100111111001110001101;
		8'd165: 64'b1101111011000101100111111001101100101111110011011100111111011011;
		8'd166: 64'b1001010110111111111111111111111011111111101111111011111111111011;
		8'd167: 64'b1110110111100011101000111100011111101101101000111000101111001011;
		8'd168: 64'b0011111001101000110111001100110110111111001110111001110111011101;
		8'd169: 64'b1101111110001111110111111111010111011110100110011100101111011111;
		8'd170: 64'b0100111100001111101110101110101100011110110011100000101101001010;
		8'd171: 64'b0111110111101100001011101010011101111111011011010000110010001001;
		8'd172: 64'b1110111110111111001010111111100101101011110111111011110001110011;
		8'd173: 64'b0011011111000011000000111100101011001101111000101101001110011110;
		8'd174: 64'b1011111111100111111111101111110001111100100111010111111010111001;
		8'd175: 64'b1011011011111011101110111111101110111010111110111111100011111011;
		8'd176: 64'b0111111100111111011111111111101101110101111111010111111111111111;
		8'd177: 64'b0011101011011111101111000111110010111000101101001011100111110101;
		8'd178: 64'b0011111111110011101001100001100011110101000001100011010100000011;
		8'd179: 64'b1111111011100111111111111011011111111111111001101110011011110110;
		8'd180: 64'b1011001100100010101110010000111110111010010111011101010001100011;
		8'd181: 64'b1101000111110010011110101110011011011001001011100111110011110110;
		8'd182: 64'b1100111011111010110010111101111010101011111110100010100110001100;
		8'd183: 64'b0111010010111001001111011010110100111011111111111111011111001101;
		8'd184: 64'b0110100110101111001111101100011101101111000001111111111111010000;
		8'd185: 64'b1101010101011101111010101110101101011100010111111101100111001101;
		8'd186: 64'b1101001101110111111010001101101111011000011101000110100101111011;
		8'd187: 64'b1101010101101011001111010001100111111101011001110011111110001111;
		8'd188: 64'b0111111010001010010111011101110010011100110011100001111001011101;
		8'd189: 64'b0110101010010111101100010110011101100001010110111100010110101110;
		8'd190: 64'b0001110111110010110101110110010111011111001111111111011011100111;
		8'd191: 64'b1100101001111110111011100001101100111011010110101111111100111011;
		8'd192: 64'b1110011101111111111111111111101111100111011011111101011101101000;
		8'd193: 64'b0111010001101101011101111000111101111111100010110011111101000111;
		8'd194: 64'b1111011101111101110110111111011111010111111101011101011101011101;
		8'd195: 64'b1100101000010111110111010011111010000001100101011001110101111101;
		8'd196: 64'b1111000110011001010100010000110001000110110110100101011110111100;
		8'd197: 64'b1011011111100010101101111011101011101111101111101011101100111011;
		8'd198: 64'b0010101010111111110001110010110101100011110111111111110111111101;
		8'd199: 64'b0111111111001111011001001110111111110110110011100101010111100011;
		8'd200: 64'b1101011110110001111111110011100000011100110100101101110010111110;
		8'd201: 64'b1101001001110011111100001011000110110001000100111111111000100011;
		8'd202: 64'b1011100110101110011010110010101000101000111101111111101000110011;
		8'd203: 64'b0110011010101110100101110100111001101111100001100011011111111111;
		8'd204: 64'b1111110010111110100110111010010111101110111111101101001010001110;
		8'd205: 64'b0100011010110101111110110000000110011100011001111011000010011100;
		8'd206: 64'b0111101110101001111111101011010101111000101010010110110110110000;
		8'd207: 64'b0110111111101011101101110110001111101110110011111011011101011010;
		8'd208: 64'b1001101111101011101101111011101111111011010110111011110001000011;
		8'd209: 64'b1111001111111110101110110111010111010001011111110000010101010101;
		8'd210: 64'b1111110100111111111011010111111111111010111111111000101111111111;
		8'd211: 64'b1111011011111111101111101011111111111110011111110101110110111111;
		8'd212: 64'b1000011101000010110101111110111010100111101010111100001101000111;
		8'd213: 64'b0001111000111111101011111011011100010110111111111010111001111111;
		8'd214: 64'b1101100100111111011110011111001100110100000100110111010010111010;
		8'd215: 64'b1110111111100111101111111011111101101111111100111101111011101011;
		8'd216: 64'b1111011011111010100111010111101011111010001111101111010101111111;
		8'd217: 64'b1101100100111111111101111111111011110101001111111111011000011110;
		8'd218: 64'b0111011010110111100111100111011101111011001111111111011001000111;
		8'd219: 64'b0111100101111001010111000111101100101101110011011100110001011011;
		8'd220: 64'b1011000101011100001100101011111110100000010111000111100010011001;
		8'd221: 64'b1011000111101101001110011101101010110111011110010011000011100111;
		8'd222: 64'b1110101101111011101111111111111101101011110111111111001011000011;
		8'd223: 64'b0001111111111110111110111000010010001111100110011011110010000110;
		8'd224: 64'b1011111111111011101101101110101010110111011010011111111111101011;
		8'd225: 64'b0110011010011100101110101000110011100001101000100010111010010101;
		8'd226: 64'b1110111111111111111011011101011101001110011110111101110101101110;
		8'd227: 64'b1110111001010110110111011100111111001100110111100100111111101111;
		8'd228: 64'b1011101110011100000110111001111010011001110110000010000111011001;
		8'd229: 64'b0011011010100100011111101000000100100001011011001110111001010000;
		8'd230: 64'b0001001111011011011110010001011110110011000111111000001110111011;
		8'd231: 64'b1111101101111110101011111011110111111010011010100010111010101111;
		8'd232: 64'b1111111111111111111011101111110111111111111011111111111011101100;
		8'd233: 64'b1010110110101001110010011010001110011011111011001010011110101000;
		8'd234: 64'b1011111011110101011111001101100110110111110100011101111011011010;
		8'd235: 64'b0111110101000001111110100111010010011011011001100101100001100010;
		8'd236: 64'b0100100111011001010111110011000011111101101101101100110101111011;
		8'd237: 64'b0100110101101110011011101111011111111111011011110101010111101100;
		8'd238: 64'b0110010111011111101110000101011110111011110000111110111011101001;
		8'd239: 64'b1010111011111100111111111101110110001101110010111001111101111101;
		8'd240: 64'b0111011101110101010101110111011011111001010100111101110100111001;
		8'd241: 64'b1111001111111111110011101111110111010111110111110101101010011111;
		8'd242: 64'b0010000111111111010100000011101000100010001011110001010011111010;
		8'd243: 64'b0101111011101011110001100110001100111011001011101111011000101111;
		8'd244: 64'b1110101101011101111110001111010101100111111111011111011111111110;
		8'd245: 64'b1010110111111000100001001100100011100101111111110000010010011110;
		8'd246: 64'b1101110101000011011101011011101011110100010101011101000101011111;
		8'd247: 64'b1011111110110110111101110011110110011111111111010110101111011001;
		8'd248: 64'b0110111001111011111010000111111111100111000100111110111101111100;
		8'd249: 64'b1111110100110011010011101111101010000101101100100101001100011011;
		8'd250: 64'b0100100000001011000111111100101000110101111010010001110011001010;
		8'd251: 64'b1100011011100111110101100110110111100101111001000101111000110110;
		8'd252: 64'b1101100111100110111110000010100111101101000101101111101001101101;
		8'd253: 64'b1101101101101111101101000111111111010111011111110011111110111111;
		8'd254: 64'b1001111010111101111111111110101111111101111111101101111011001110;
		8'd255: 64'b1001000111101010111110011100101110101011111101011110110111011010;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page6(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1101011101111001101111100111010111010100111101001011010101110111;
		8'd1: 64'b1101011111100111111111101111111111110110111101110110111110111111;
		8'd2: 64'b1111111110010110001011111101001110110111100101100010111111111111;
		8'd3: 64'b1101111000111000111111001011011110011100000100001010010101010011;
		8'd4: 64'b1111000011110110010100011111101111110000111011010111011101111100;
		8'd5: 64'b0111111011111101111001111111010111111111111011011111111111111101;
		8'd6: 64'b1111101101101011110011110001100001111001111110101110101101111000;
		8'd7: 64'b0000011101010001010011000000110010101111001011100010000110000000;
		8'd8: 64'b1011111111111111101100010001000100111001001111100011101100011111;
		8'd9: 64'b1110101111111010001011110000111110111011100111101010111100010111;
		8'd10: 64'b0110001101111011110101101111101011000110111110101111111011111010;
		8'd11: 64'b1111100111011110010010001110101111001101111011110111111111111111;
		8'd12: 64'b1100111111111010100111101011011101011111110111101101111011111111;
		8'd13: 64'b1111101111000111010111001100010011011110000100001101101101000001;
		8'd14: 64'b0001011110111110000111110110011111010111110101100011010100111111;
		8'd15: 64'b1111010011000101111011001010010001111110101111011111110101111111;
		8'd16: 64'b1111100111111100101001011111110111101011110011111110111001011011;
		8'd17: 64'b0101101110101101011010101100100110101101111011111100001010100101;
		8'd18: 64'b1101111110110111011110111110111101110111100101101111111100101110;
		8'd19: 64'b0111100100010011111101111011001111011001011011111101011101111111;
		8'd20: 64'b1110100110111000111111101110101111001101101011101011111011101010;
		8'd21: 64'b1001101011100010101011111110001110111111110000111010111011111111;
		8'd22: 64'b1111101011110111110011001010101111000100111111101111110110111011;
		8'd23: 64'b0110001010111101110111100111111101101111101110111110111101111111;
		8'd24: 64'b1111111000001110111111011010100111101100111111001111111011100111;
		8'd25: 64'b0111101110101011111111111011011111101010000101010011101010100010;
		8'd26: 64'b0111010001001101111100111100010011011010111011001100101111101101;
		8'd27: 64'b1100111111011111111111111101011011101011111101111110111111011100;
		8'd28: 64'b1110111010101110101111111111111101111110101011110110111011111110;
		8'd29: 64'b1011100111010111100011110010011110011111110001001011111101101001;
		8'd30: 64'b0101111110010010010001110101001001101011011001100101001111001010;
		8'd31: 64'b0111100100010110110101011101100111110001000010011100111011101011;
		8'd32: 64'b1111111111101011000110111101100011111111111001111110101111011101;
		8'd33: 64'b1111111011011111111111010100011111111110100101011110110100110101;
		8'd34: 64'b0111111110101111100011111111011011110111100101110111011111100111;
		8'd35: 64'b0100110101000011010100111010101111001111110111010001001100111100;
		8'd36: 64'b1100010001000101101000111111111100011111010011111111101111001101;
		8'd37: 64'b0110101001100100111110011111001011111000101011010011111111110000;
		8'd38: 64'b1111111101111011100001110100001011001111111101011101011111000011;
		8'd39: 64'b1011001011111110110101011011110111110111111111111111011100011101;
		8'd40: 64'b0101111111001111000001101111101111111110111001111010011111111111;
		8'd41: 64'b1101101100010110000110100111101100001110110011101010101100011110;
		8'd42: 64'b1100101111111100011110111110101010111000011110100110011101101001;
		8'd43: 64'b1011111111001101111111110111010110011111101111111011011010110100;
		8'd44: 64'b1100011001010101000111111101101111001010011010011111111111011011;
		8'd45: 64'b0111111101010110110111010001111101110111010011111101110010111011;
		8'd46: 64'b1000110000111001101011011101111110001100001111001001111101001111;
		8'd47: 64'b0111011101110010101000101111001101110101011111000010011000001000;
		8'd48: 64'b1111011111101001101010110110010110101111010111111111100101111101;
		8'd49: 64'b1111100101111101110111111111000100111010011110111001111110111111;
		8'd50: 64'b0001111011011001111111111111111111111110110011011111111011111111;
		8'd51: 64'b1111111110000110101001100111111111110011111000110110111110111000;
		8'd52: 64'b1101110001011001111111110100100101111011111001010101100001011011;
		8'd53: 64'b1111100011110101011111110101011111111001011101111011110111111111;
		8'd54: 64'b1000111110110110111001100111111000100110000111101010111011111110;
		8'd55: 64'b1010111111101110110110111111101110011000101110111111011111110111;
		8'd56: 64'b1100011001011100101011001000011010001010011011011110010011001010;
		8'd57: 64'b1101100111111101011000111101000111011011011110011110010101100111;
		8'd58: 64'b1101000111110111110110001111101011010101010101101101100101111110;
		8'd59: 64'b0010111001111001101001110110001001100110011111010011111101110010;
		8'd60: 64'b1111111000111111111111111111111110011100011011100111111011111111;
		8'd61: 64'b0110101010111101111011001011100111111111111011110010110111011111;
		8'd62: 64'b1110111011101000111111011101101111100110111011011011011111011111;
		8'd63: 64'b1011100010001101110110001011111101111110101110100001111101001011;
		8'd64: 64'b1111111101111011001001110011001110111111111101110011011111110111;
		8'd65: 64'b0011100010010111111110000011100010111110111101001111000111111110;
		8'd66: 64'b1111101011011111101111001101111111111100111111111010000111011101;
		8'd67: 64'b0011111000110001000011111011110010111011111100001010111111111111;
		8'd68: 64'b1010010011101101001001001000111010000100111011111110010110001000;
		8'd69: 64'b1111101101001011100100000111101100011111101010111001100000011010;
		8'd70: 64'b1001110110110100000010101111111010011000010111111000100011111110;
		8'd71: 64'b0010110111001110000001111001111000101110011011000010111010011110;
		8'd72: 64'b1110011111111111111110111101101000101111111001111010101111100110;
		8'd73: 64'b1111101010000100011111001110010111111111111111110101101001100111;
		8'd74: 64'b0111111111110111011011111110011111111111011100111101111111111101;
		8'd75: 64'b1101100111001011111011110001101100101001000110101000111101001111;
		8'd76: 64'b1101110011011110111111101101111111011110111101111111110011110111;
		8'd77: 64'b1111111011010011110001111111111111111101110100111100100111100111;
		8'd78: 64'b1111110111011100111011101101111011101100110111001111110001011101;
		8'd79: 64'b1110011110101001111111110001101100100101001111111111010100010001;
		8'd80: 64'b1111011111110101111111100111011111110111011101100111011100110110;
		8'd81: 64'b1100011111111011010001111110110101001111111010111110111110101101;
		8'd82: 64'b1111100111100101111111011101011010110111110001101101110111010000;
		8'd83: 64'b1110101110101111111011110000110011111100111010111110111110101110;
		8'd84: 64'b0110111111101111111111110011111101100101011111010100101110011100;
		8'd85: 64'b0011111101100111001100100110011101101110111111110010111111100110;
		8'd86: 64'b1110111101001110001111100110111100111111010001011111111111101111;
		8'd87: 64'b1111100011101110111001011110110100101110011011101010100010001011;
		8'd88: 64'b1010001111101110111110110011111010100110111111111111111110011110;
		8'd89: 64'b1101110010110000110100110101110000011100111100011110011111111100;
		8'd90: 64'b1101010110110111000011111101110111011011101110101110111111010100;
		8'd91: 64'b0011110101110001111001010011101011111111110000000101110000110110;
		8'd92: 64'b0111110111100111111011001101000101111101010100011011100011011011;
		8'd93: 64'b1010111110101000101011101010100110101101111010001101101101001011;
		8'd94: 64'b1101101111111111110111111111101001011111111111101001101101000110;
		8'd95: 64'b1111010110001111010001010111111001010110111011010111111010011011;
		8'd96: 64'b1011111101111010100111111001001011111011110111111001111111110111;
		8'd97: 64'b1010111111111111110111110101011111101111001001001001111100100111;
		8'd98: 64'b1110010111111011011101111111111101110111111110111101111101101011;
		8'd99: 64'b1011111001110010111011100111111010110111111101000110001101110010;
		8'd100: 64'b1001101111001101100111101010111010011001101011001111111110101111;
		8'd101: 64'b1110110110111111111111101110011111010010101011111011011010001111;
		8'd102: 64'b0011101010011111011110100011010011111110110111100111111110001000;
		8'd103: 64'b1111010111110110111110100101001111111111110101000111111101110110;
		8'd104: 64'b1111111101000111010111110001101110110011101101111111101111011011;
		8'd105: 64'b1111111111101101011110111110110011101111110111010101111110000100;
		8'd106: 64'b0100101101111011010001100100101011111011111111110100001101011110;
		8'd107: 64'b1101010101010111010010100010111111011100100111000110001101011110;
		8'd108: 64'b1010101011101100011001101010101011110110101111101110011110111010;
		8'd109: 64'b1110010100001101110010011010011110010111001110010111100111110111;
		8'd110: 64'b0101110011101111000100101011111011011011111101101111111001110100;
		8'd111: 64'b1101101111011111110110010110011101110101100100111111101100110111;
		8'd112: 64'b1011011110011101110111110010011111011111011110111111111101101111;
		8'd113: 64'b1001100000011011101100001111101111011100000111111011010001010111;
		8'd114: 64'b1011110010101101101011001001110111101111111111010001110110111001;
		8'd115: 64'b0100010110111111011111011100101011110101011110100111010000101110;
		8'd116: 64'b0110011100111111001010011101011110110111001100111111111001111110;
		8'd117: 64'b0111011111111111001110100111001101100111111011110110111111111111;
		8'd118: 64'b1111111111001011110000011011111011011010111111111110001111101111;
		8'd119: 64'b1100111010110110100111111001001011111110110111111001111110011111;
		8'd120: 64'b1100101110110111011010101101111100111011111101110110111110100011;
		8'd121: 64'b0111111111111100111010100111101011110100111110001110001111100000;
		8'd122: 64'b0110111100100111011111100010111101110110111001110110101111100110;
		8'd123: 64'b0110000111100111111110011111111011100000011110111110000101101111;
		8'd124: 64'b0101100000110011100001011011111101010001111100101010000111111110;
		8'd125: 64'b0111101101011011101111110001010111111000111101110011010101110011;
		8'd126: 64'b1011001100111110100111101110111011000111111011101110101110001111;
		8'd127: 64'b1011111101101111111011110110011100110111011001010010011100101101;
		8'd128: 64'b1001110110111110101111111100101111111000110111101111111011011011;
		8'd129: 64'b1001110111011111110111011111010111111001101111010010001111100000;
		8'd130: 64'b1101010111111101110100000101111110011111111111011101011101011111;
		8'd131: 64'b1101110111010001111111011010100011101011111000111111111011101000;
		8'd132: 64'b0111111111111111101110111011111101110101100100111111111110001111;
		8'd133: 64'b1001111110111101101011111101101111011011011111011111111001011011;
		8'd134: 64'b0100110111001011110011111111100111111111111011101110111111011000;
		8'd135: 64'b0111011101111011000011100111101000111111111100110110111111111010;
		8'd136: 64'b1110011011011101100001111110101011101111111011011010111111001110;
		8'd137: 64'b1101011111110101101101111111111110010001111111111001000111110101;
		8'd138: 64'b0111010111010111111101111101111111111111010111110111010001101100;
		8'd139: 64'b0101110010111011111011111111100110000101001111101111100101110111;
		8'd140: 64'b0000101011001100110011011000010101001010110101100000111011011000;
		8'd141: 64'b0100100110111110001110111010111110010110101101000010111110111101;
		8'd142: 64'b1110111110111111111111000111111111101110101111111110111011111101;
		8'd143: 64'b1110111111101011000101111110011100111011001111110111001101101111;
		8'd144: 64'b1011010111111101101100011111100010111101101111111001111010111100;
		8'd145: 64'b0111111111111101011001011101111110110110111011100100011101111111;
		8'd146: 64'b1110110111111110111010011110110010101111111111101010110111111101;
		8'd147: 64'b0110111001000101110110111011101111110011101000111101110010010010;
		8'd148: 64'b1100011110000111110100011001110011001000101010100001101000100100;
		8'd149: 64'b1011101101110110100011111111011110111011011111100000101001101110;
		8'd150: 64'b1111110110110111111111011011011111101001111101110111111111110111;
		8'd151: 64'b1101010101110011101111000101101010110110011110011011010111000100;
		8'd152: 64'b1111111011101111111011111111111111111110111111111110111111111111;
		8'd153: 64'b1111111110010011101111111001111111111011101110011111111110111011;
		8'd154: 64'b0110110101101011111011111111001101001111111011111110111111001110;
		8'd155: 64'b1100111100110110110111010010110011111100110001110101110001110110;
		8'd156: 64'b1111101111111111111011110101001111011001011111110111111100111010;
		8'd157: 64'b0111010111011000110100011111110011010011110010001101000111111011;
		8'd158: 64'b0110110111011111011101101110011101101101101011011100010011110111;
		8'd159: 64'b1011110111110110101100101111101010110000011011110011011111111110;
		8'd160: 64'b0111110100010111101001111111110101110111111011010100011101001101;
		8'd161: 64'b1010101010110110111111111011101010111101001111101110010110111010;
		8'd162: 64'b1111111011011011111111011101101001101110110110100100100111111011;
		8'd163: 64'b1111011111111011111101101111101011111111111110111101011011111010;
		8'd164: 64'b1001100100011101000111010011111110001011100100111111001110001101;
		8'd165: 64'b1101111011000101100111111101101100101111110011011100111111011011;
		8'd166: 64'b1001010110111111111111111111111011111111101111111111111111111011;
		8'd167: 64'b1110110111100011101010111100011111101101101100111001101111001011;
		8'd168: 64'b0011111001101000110111011101110110111111001110111101110111011101;
		8'd169: 64'b1101111111001111110111111111110111011110100110011100111111011111;
		8'd170: 64'b0100111100001111101110101110101100011110110011100000101101001010;
		8'd171: 64'b0111111111101100001011101010011101111111011111010000110010011101;
		8'd172: 64'b1110111110111111001010111111100101101011110111111011110101110011;
		8'd173: 64'b0011011111001011000000111100101011011101111000101101001110011110;
		8'd174: 64'b1011111111100111111111101111110011111101100111110111111010111001;
		8'd175: 64'b1111111011111011101110111111101110111010111110111111100011111011;
		8'd176: 64'b0111111100111111011111111111111101110101111111010111111111111111;
		8'd177: 64'b0111101111011111101111011111110010111000101101001011100111110101;
		8'd178: 64'b0011111111110011101001100001100011110101000001100011010100000011;
		8'd179: 64'b1111111011100111111111111111011111111111111001101110011011110110;
		8'd180: 64'b1011001100101010101110010000111110111110010111011101110001100011;
		8'd181: 64'b1101000111110010011110101110011011011001111111100111111011110110;
		8'd182: 64'b1100111111111010110010111101111010101011111110101011100110001100;
		8'd183: 64'b0111110110111001101111011011110100111111111111111111011111001101;
		8'd184: 64'b0110100110101111101111101101011101101111001001111111111111011100;
		8'd185: 64'b1101010101011101111010101111101101011100110111111101100111001101;
		8'd186: 64'b1101001101110111111010001101101111011000011101010110100101111011;
		8'd187: 64'b1111010101101011001111010001100111111101011001110011111110001111;
		8'd188: 64'b0111111010001010010111011101110010011101110011100001111001011101;
		8'd189: 64'b0110101010010111101100011110011101100011010110111100010110101110;
		8'd190: 64'b0001110111110010110101110111010111011111001111111111011011100111;
		8'd191: 64'b1100101001111110111011100011101100111111010110111111111100111011;
		8'd192: 64'b1111011101111111111111111111101111100111011011111101011101111000;
		8'd193: 64'b0111011001101111011101111000111111111111100010110011111101000111;
		8'd194: 64'b1111111101111101110110111111011111010111111111011101011101011101;
		8'd195: 64'b1100101000010111110111010011111010000001100111011001110101111101;
		8'd196: 64'b1111000110011001010100111000110001000110110110100101011110111100;
		8'd197: 64'b1011011111100010101101111011101011101111101111101011101100111011;
		8'd198: 64'b0010101010111111110001110010111101100011110111111111110111111101;
		8'd199: 64'b0111111111001111011001001110111111110110111011100101011111100111;
		8'd200: 64'b1101011110110001111111110011100000011100110100101101110010111110;
		8'd201: 64'b1101011101110011111100001011001110110001000100111111111000100011;
		8'd202: 64'b1111101110101110011010110010101000101000111101111111101000110011;
		8'd203: 64'b0111011010101110100101111100111001101111100001100011011111111111;
		8'd204: 64'b1111110010111110100110111010010111101110111111101101001010001110;
		8'd205: 64'b0100011010110101111110110001000110011100011001111011000010011100;
		8'd206: 64'b0111101110101001111111101011010101111000101010010110110110111001;
		8'd207: 64'b0110111111101011101101110110001111111111110011111011011101011010;
		8'd208: 64'b1101101111101011101101111011101111111011010110111011111001001011;
		8'd209: 64'b1111101111111110101110110111010111010001011111110001010101010101;
		8'd210: 64'b1111110101111111111011010111111111111010111111111001101111111111;
		8'd211: 64'b1111011011111111101111101011111111111110011111110111110110111111;
		8'd212: 64'b1000011101010010110101111110111010100111111010111100001111100111;
		8'd213: 64'b1001111000111111101011111011111100010110111111111010111001111111;
		8'd214: 64'b1101100100111111011110011111001100110100000100110111010010111011;
		8'd215: 64'b1110111111100111101111111011111101101111111100111101111011101011;
		8'd216: 64'b1111011011111010100111110111101011111110001111101111010101111111;
		8'd217: 64'b1101110100111111111101111111111011110101001111111111011100011110;
		8'd218: 64'b0111011010110111100111100111011101111011001111111111111001000111;
		8'd219: 64'b0111100111111001010111000111101100101101110011011100110001011011;
		8'd220: 64'b1011000101011100001110101011111110100000010111011111100010011001;
		8'd221: 64'b1011000111101111001110011101101110110111011110010011000111110111;
		8'd222: 64'b1110101101111011101111111111111101101011110111111111001011000011;
		8'd223: 64'b0001111111111110111110111010010010001111101110011011111010000110;
		8'd224: 64'b1011111111111011101101101110101010110111011010011111111111101011;
		8'd225: 64'b0111011010011100101110101000110011100001101000100110111010010101;
		8'd226: 64'b1110111111111111111011011101011101001110011111111101110101101110;
		8'd227: 64'b1110111001010110110111011100111111001100110111100100111111111111;
		8'd228: 64'b1011101110011100000110111001111010011011110110000010100111011001;
		8'd229: 64'b0011011010100100011111101000000100100001011011001110111001010000;
		8'd230: 64'b1011011111011011011110010011011110110011000111111000001110111011;
		8'd231: 64'b1111101101111110101011111011111111111010111011100010111011101111;
		8'd232: 64'b1111111111111111111111101111110111111111111011111111111111101101;
		8'd233: 64'b1110110110101001110010011010101110011011111011101010011110101000;
		8'd234: 64'b1011111011110101011111001101100110110111110101011101111011011011;
		8'd235: 64'b0111110101000001111110100111010011011011011001100101100001100010;
		8'd236: 64'b0100100111011101010111110011101111111101101101101100110101111011;
		8'd237: 64'b0100110101101110011011101111011111111111011011110111110111101110;
		8'd238: 64'b0111010111011111101111000101011110111011110000111111111111101001;
		8'd239: 64'b1010111011111100111111111101110110001101110110111001111101111101;
		8'd240: 64'b0111011101110101010101110111011011111001010100111101110100111101;
		8'd241: 64'b1111001111111111110011101111111111010111111111111111101010011111;
		8'd242: 64'b1010000111111111010100000011101000100010101011110001010011111110;
		8'd243: 64'b0101111011101011110001100110001100111011001011101111011000101111;
		8'd244: 64'b1110101101111101111110001111010101100111111111011111011111111110;
		8'd245: 64'b1010110111111010100001001100100011100101111111110000010010011110;
		8'd246: 64'b1101110101110011011101011011101011110100010101011101000101011111;
		8'd247: 64'b1111111111110110111101110011110110111111111111110110101111011001;
		8'd248: 64'b1110111001111011111010000111111111100111000111111110111101111100;
		8'd249: 64'b1111110100110011010011101111101010000101101100100101001100011011;
		8'd250: 64'b0100100000001011000111111100111000110101111010010001110011001010;
		8'd251: 64'b1100011011100111110101100110110111100101111001000101111000110110;
		8'd252: 64'b1101100111100110111110000010100111101101000101101111101001101101;
		8'd253: 64'b1101101101101111101101010111111111010111011111110011111110111111;
		8'd254: 64'b1001111010111101111111111110111111111101111111101101111011001110;
		8'd255: 64'b1101000111101010111110011100111110101011111101111110111111011010;
	endcase;
	return out;
endfunction
