function Bit#(256) get_msg_bit(UInt#(6) counter, UInt#(3) page_num);
	Bit#(256) msg_bit = case (page_num)
		3'd0: get_msg_bit_page0(truncate(counter));
		3'd1: get_msg_bit_page1(truncate(counter));
		3'd2: get_msg_bit_page2(truncate(counter));
		3'd3: get_msg_bit_page3(truncate(counter));
		3'd4: get_msg_bit_page4(truncate(counter));
		3'd5: get_msg_bit_page5(truncate(counter));
		3'd6: get_msg_bit_page6(truncate(counter));
	endcase;
	return msg_bit;
endfunction

function Bit#(64) get_prev_enc_page(UInt#(8) counter, UInt#(3) page_num);
	Bit#(64) prev_enc_page = case (page_num)
		3'd0: get_prev_enc_page0(counter);
		3'd1: get_prev_enc_page1(counter);
		3'd2: get_prev_enc_page2(counter);
		3'd3: get_prev_enc_page3(counter);
		3'd4: get_prev_enc_page4(counter);
		3'd5: get_prev_enc_page5(counter);
		3'd6: get_prev_enc_page6(counter);
	endcase;
	return prev_enc_page;
endfunction

function Bit#(256) get_msg_bit_page0(UInt#(5) counter);
	Bit#(256) out = case(counter)
		5'd0: 256'b0110000111110101100111001000001001111101000011100101111000010101011110001011100100011111100111010101101001100010010000010010101011101100000111001101000101111011110100000010101011101001100001100100000111010111101010001011110001011010000100111010111110111001;
		5'd1: 256'b0001101100001000101111010111001111100001001000101110101111011000101111101110000100100000001100111011001011101011111000010001000000101001101010011111001011000110100100000010110110110100100000000110010001011101100101111010101011011001010100001101100000000111;
		5'd2: 256'b0000000101010000010000010011010110100001011000010000001111101010010001001100100100011111110101110110100011011011000111110000001011111000001100011101010100010011000100000011000110000101001100010110101111101110011011000100000101100000100101011001011000001100;
		5'd3: 256'b0101100100011101010001000010101110110110111110000011111100101001111110010000011100000111000101111101001010100001110100110101101001111101100010101101111001000001000010001101100011100011000010110111011100101011100110110011001011111110100001000110000101111001;
		5'd4: 256'b0010001111110000001011001001001011101010110001000010010011100010011011000100100100111100101110100101100010110011010111101100010001010011010100000101111100000010001000001100001101001100100111110111000010101000010110101010010001001110010001100000001110010001;
		5'd5: 256'b0110011100001100010010010011111110101010101100000111010110101111010001011000011110011111101010111100100110010110101100000001001001110001100010000100011111001010110010010110000101100101010011100010100001100100100010001101001010001101100000101111010110100001;
		5'd6: 256'b1000100111100011000111010011010111001100001101100010101110101010001010100011000101010101010001100011100110101001001110110111111000100111011110101110000001001110010001000000010010110101011011111110000010001100001000110011011110001001101101001001100100100111;
		5'd7: 256'b0001100010010100101110001100001010010001111101010100110001100010010111101110010110101010111001010101111001011100111100111000010010100010101010110000010000101101010000111101001010010010000011100001100111110100100101011001111111100011001011001001001011101101;
		5'd8: 256'b1010111010001011010011001000000100000001010101100001001000011100000000000001011101101100100100111111010111110100010110100111110110000100110111011111100101011001111000111100001110001011111001101000001000101011110100100001110001111000111010111110000101111001;
		5'd9: 256'b0100110011110011000111101111001111001010111010101101001110101011111001010110100101000111001110100101001111001111101111001101111100100101110111010101110001101100110010111011100110101000010100111111011110111111011100101011000100001001111101111101111111110010;
		5'd10: 256'b0000010101000000110000001100010111100111111100000000010100011001101111110110010010000001001110001100001100100100000000000110110101111110110011111111110010111100011011000110010001010011000010001110010110000011010010101001101101101100110101100001011001001010;
		5'd11: 256'b0011011110001101110010110100100011111110001111001000000011000001101011100100011001010111111001000111000100010000101000010111000100101100110100111100010010001101010011111010110001111111110001101011100111001001011011111001110010011110101011010000000001100100;
		5'd12: 256'b1011110101110011111011110111110000101001010101010001111110001001010111010111011010101000101101100000000010001111100001100001010100001001000010000110101101110010110101010010000001101000111011000101010010111000100100101111001010010111001001011000100111011110;
		5'd13: 256'b0110000100100110101101010000111101000101100101001110101011000011101010100111010011111011001111110001110111101011001101110100011111000110101110110101000001111010000101101101110100111111011110110001101001110101001111010011000001011011101111100010110111000001;
		5'd14: 256'b1000001111100100101000010111000111100011110100100100100110110101011100110100110011101001111000010100001110100011100101001010100000100100000000011100110110111010000111111110011100110101010000111000111111100100011010100110000011011111010011001111001100010010;
		5'd15: 256'b1101100010001111001010100110011011010011011010111110110001010101101000000011011101111100100000001111011110000001001100110000001101100101001000101110011000000100011011101010000100100101101010100110101110011000000011111101100110000101000100110011011000010111;
		5'd16: 256'b1110110001110001000000110011101101000111001010011110011011101111101001111100110110011001100000010110101000111110000101101011010010001111111111110100100110110111100000101000111111101010010110001001100001010000110111101000001011001011100100000100011000101100;
		5'd17: 256'b1010011101001110010100011101011001010110100101010011110110010110111000010110110011110100000011001011011010011001111111111110101010101001101101000011110111110011100001111110100000000100001001010111011011101001100011110101001111010001111110101100011101000011;
		5'd18: 256'b1010010000101110001000001101001001110010011001000101000001000101110101101101101000011111101110101011000011101000111100100110001101100001101110111001001011101111000111001110001110010110111101010011100111001001111111100000000000111001010111000001001000101101;
		5'd19: 256'b1001011011011000110011100001100111111010010011001101111101010101011000110011011110000000100100001010110010001100101000001111110110011100100100111110000100110000000110101001100110010111011110001100000001111101111111000111000001000000111110111110011011001110;
		5'd20: 256'b1000001001110101000001010111010011101100001111001110010010100010001001101101110111000100100100101000011110001000000101101001100001000100011101001011000010111111101101101010010010111000010010001110111001101011001110111000011101110011000011110011011010010011;
		5'd21: 256'b1100101111010010001101101101111001100100110010110011011011001110101111001010111101111101000010101111100011001100011011110010001101001011010101010010011111001010000011111101000101011001101101001101101111110000101001010000111101111110010110110110110100011100;
		5'd22: 256'b0000100010100000000101111011110010011010110101001001101010101100100001111010011000001101001111000010110001001100011111100000100001100011011111011010111001110000101001101010011001000110011001100100101000001100011010000010010111011110100010111001111010011111;
		5'd23: 256'b1110011100111110010100101101001010010011001011000110001001101001111110101101110101010111111010100011111000010110001110000110110110010101101010011110110110100010111011101100001000110110011101010101101110101010001001111111000000011010011110100011010101110101;
		5'd24: 256'b1001111010100010010000001011001011001111010110010011110000111010010010110000010111001000001100001011101010101110001011011011011001111101110010010100001110000100101100010001001101100010010110101010111000100010110000011111011001110001011001001000100110110011;
		5'd25: 256'b0110100000110101101110110100110010011110011110001011001110000011101001001011010001101111011101110110100001111100001111011110110110000011011011100110010100011101010110000101101000111010001110111000001111011110101011100110101011010110001000001000111111100100;
		5'd26: 256'b0000011010101101010011101001001101010010101110110011000010010111000111001101010110111110000111111101111010110000110010111001110110011000001000101000010001010110100110001010101101001111010110011100000110110000001000011010111111001100010101001101111011111000;
		5'd27: 256'b0100001000000011001111011011101011110000101101001001101110110011110111001011110000111101110001010010101010100001000001101100001111001111001010100001010000010011100111110100110110001111011011011001001000001000001101011110110111000110000001110001100110101000;
		5'd28: 256'b0101011110111101100111100001101100111111111000100000110010111100101000011111111001010100001110011010111010001100010010110010111101100000101100101101101000011001010000101111110010000010000110101000100001110100001101011010111001100010011001101101100101010010;
		5'd29: 256'b0001110010010111001101110110011100101010001110011011101011100110101101101001001010111101101000001011011001011001011011101110001011011010101100000100110001100000110010011111101010111100111000001010010010000010001111011100100101000000100110001111111100100011;
		5'd30: 256'b0110011001000000010011110110000010010111110111110011101101010101001000000010111111011000001110100101001101000000101000011111011000110100110110111111111111110111100000110100101111000011111101000010101000101100000100010100101101001010011110110010010010100111;
		5'd31: 256'b1111111001101010100110000101001111110000101010011111000000011110010010000000111010011011111001011011001110100101010101111110000110001111111100110100000011011011101011000101000111011010100010001101001100110100010010010100101101011011110100110000001100000111;
	endcase;
	return out;
endfunction
function Bit#(64) get_prev_enc_page0(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd1: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd2: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd3: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd4: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd5: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd6: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd7: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd8: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd9: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd10: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd11: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd12: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd13: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd14: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd15: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd16: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd17: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd18: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd19: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd20: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd21: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd22: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd23: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd24: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd25: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd26: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd27: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd28: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd29: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd30: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd31: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd32: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd33: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd34: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd35: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd36: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd37: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd38: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd39: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd40: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd41: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd42: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd43: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd44: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd45: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd46: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd47: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd48: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd49: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd50: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd51: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd52: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd53: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd54: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd55: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd56: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd57: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd58: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd59: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd60: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd61: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd62: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd63: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd64: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd65: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd66: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd67: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd68: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd69: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd70: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd71: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd72: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd73: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd74: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd75: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd76: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd77: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd78: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd79: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd80: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd81: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd82: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd83: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd84: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd85: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd86: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd87: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd88: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd89: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd90: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd91: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd92: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd93: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd94: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd95: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd96: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd97: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd98: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd99: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd100: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd101: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd102: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd103: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd104: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd105: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd106: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd107: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd108: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd109: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd110: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd111: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd112: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd113: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd114: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd115: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd116: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd117: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd118: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd119: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd120: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd121: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd122: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd123: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd124: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd125: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd126: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd127: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd128: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd129: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd130: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd131: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd132: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd133: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd134: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd135: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd136: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd137: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd138: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd139: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd140: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd141: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd142: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd143: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd144: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd145: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd146: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd147: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd148: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd149: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd150: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd151: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd152: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd153: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd154: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd155: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd156: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd157: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd158: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd159: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd160: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd161: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd162: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd163: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd164: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd165: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd166: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd167: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd168: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd169: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd170: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd171: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd172: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd173: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd174: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd175: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd176: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd177: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd178: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd179: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd180: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd181: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd182: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd183: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd184: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd185: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd186: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd187: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd188: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd189: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd190: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd191: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd192: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd193: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd194: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd195: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd196: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd197: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd198: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd199: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd200: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd201: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd202: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd203: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd204: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd205: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd206: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd207: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd208: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd209: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd210: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd211: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd212: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd213: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd214: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd215: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd216: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd217: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd218: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd219: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd220: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd221: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd222: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd223: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd224: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd225: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd226: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd227: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd228: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd229: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd230: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd231: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd232: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd233: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd234: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd235: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd236: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd237: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd238: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd239: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd240: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd241: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd242: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd243: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd244: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd245: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd246: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd247: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd248: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd249: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd250: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd251: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd252: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd253: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd254: 64'b0000000000000000000000000000000000000000000000000000000000000000;
		8'd255: 64'b0000000000000000000000000000000000000000000000000000000000000000;
	endcase;
	return out;
endfunction
function Bit#(256) get_msg_bit_page1(UInt#(5) counter);
	Bit#(256) out = case(counter)
		5'd0: 256'b1111110000101110101110011100111001000100001000011111001010100100110100001100101000101100001000001011000100101000101011110100110111100100101101000110111100111100010010010111010100011011000110110110000010011011000010011011001111010111101100000010010010000010;
		5'd1: 256'b1000000111000011011111001100011101000000001101101101100001111011001110010110001110011001000001000111111100010001100010101010100110011010101011100011101010101111001101011000000000001111011110010011110000001010011111010110101010110000011100111111100101111001;
		5'd2: 256'b0011010100010001111010001111010111111111111011010010100110011101010110101000101111011011110101010011011000111000111010001010100010000100010111011100001010111011110101000110101110101001011100110111001001100101011110111100011000100101010001101011011100111000;
		5'd3: 256'b0011101101111101001101000110110111010000011011010100110111011000111100011101011010010111010001100010110100001011011000010010100111011111000000000110000111101110100001010110001101001010011010011001011111010110111110110111100000100100000001011000111100011101;
		5'd4: 256'b1000000000111110001100001101101100100100111000101001111100101000000110010011110110111100101101110110011111000001100111011100001010000110001110110100101110110000101110011110100010111000011101001010100011110101011000100010001111010010101110101101001001110001;
		5'd5: 256'b0000100010110100100111101011111111111111001011011100010001010011101011111110001110101010110010101110010111101111001001100110110000101001010011010001100101001010101011100111000011111100011011111010000011011010110101000101001101111101100001001101011100100111;
		5'd6: 256'b0000010110100101001001110111111101000110001101010011101111001000101000000101101110111101000101010111101000010010011110110001101100110000001000010110010100010011000111110011000010111001000111000000110110110110001010011000100001011101110010111001011001011100;
		5'd7: 256'b0011011011001111101101000101011111000100111111101011011100010111101111001001000010100101111110001010010101100110001011110011100101110100101111110010110011110101010111101001111010010111100111100110011010001011010110001011110011000111100110001010001111001011;
		5'd8: 256'b1100011111101100101101001100001000100100100000101010110011000100001000110010000010101010010101011000000000110000101100000111000000011100111111010001110011000101110010110001000000000011110001011100111100100001100001110011001010110000101101111111110001010001;
		5'd9: 256'b1000011111011000110010110110010101110011000001101100111110100100110111111001101111110001011010010001000110000110001011010001110001010100011000001101101011100101011100111000000010000111000001001111110111110100001101111001000011010111010110010100100011011010;
		5'd10: 256'b1101000011101010111010101110010010010001111010110011111011110010111011101011011011001101111011100111001010110111010011101101010100011010101110111101000001001001100000100110110001101101000110001001000001000101101110011100000010000111101110101000001001100001;
		5'd11: 256'b1000000000111100111111010011100011101101101101111010110111011110111101110010110000011111101010101010110111111110011000000000100110111010110100011010000110111110011110111100000001110010110110011000111010001000000001110010110110100001110110001001000110101010;
		5'd12: 256'b0111000111010010110001011010110110101110010100010011010000110110000000011011100100001001000111100100100000011101101110101100100100000111000110011101111000000110100110101100011110010101001100100110100100011111001101010110011010000111100100001011000101110100;
		5'd13: 256'b0000101001011101111010101110001011001111010101100110100000001010101000101000010011101100111111111010100011100011011001011010111000001000000111111100100100100100100001001100001111000000001001111001000100100111010010110100100101111111101101110010101001101111;
		5'd14: 256'b1110001110101110011001011101011001011111100101110100110101001110000010001000011110011110111001001110010000101101100000010111101010100111100000011101000110001000011000110011011011110000111001100011011011111111110110010101101111011100101000010110001011110111;
		5'd15: 256'b0100110010001001000111101001100110010001001011001000001010111010110100101100100001011110011000010101000001111011100001100010100011100011101010101101010110101100011101101101001001111001111110111001011100111111111011000011101000101001011101100110001001000010;
		5'd16: 256'b0100110111101000111100011011001010001011110010010011011001110111001101001100011011000011010001001110101000100111011111010011100010111011000111110101001111100010001011111001001101000000101001101001100110001101110001001010100011000110100010110110100100001110;
		5'd17: 256'b1110011100101010110101101110111101010000100011110100101011100000111000111111011110010011100101000111101101110100100001111100101110000000001101011100010011110011010100101110010001101000010010110010010011011101110100011111010111000011101100001001100000010001;
		5'd18: 256'b1010110011001011001110001101011010011110001110001010110010010010111011111000000111001100001100000110101111011100101001101110010101101110010110110101011110010100101011101010100011110011011110010100011011010000101010010110000110100011000010000000011011001110;
		5'd19: 256'b0111001001010011110000001011111010111110000010100011001100010000101110010110010101111101001110011001101111110011000001010000010111001011100011100100010000001011110101101010110001000001010001000000100010010000101110011111100011010100111101010110011000101100;
		5'd20: 256'b1101111010011111010001101101010100111011010101111011111100110001000001000111010001110101100001100011101101100100110010011101000101001110100100111001101010110101010110011000001111101010110000110000011001101100010001010101010000001000111100011010101101101010;
		5'd21: 256'b0111000000111111100111110011100011111010011100010100110001101010100010110011101101011011000000001100101011010000111000110111111001100000100101001100000100010100011111010110101011010110001000111110100010101111000011001011000010110110100110011000111001011111;
		5'd22: 256'b0000110011000100100010110011000000110101011010011010010010000001010111101111110000001101100110011011001000001101001111101100011011011110011100000001111011100111101000000111111111111011101101111100100110011101011110100100110100110000001111111110001011101101;
		5'd23: 256'b0110000110100101100101010111010101100111001011001111000100110011110000101100011101110011010000110000111110010010100111111101010110100010111111100010010100000111110000111011010100111100000110100000110111100110010110000001000010011101010111100010001000110010;
		5'd24: 256'b1000001011101001000010010000100011111101000101111000010100001001101010111110111110010100111111111111100110011101000101101011101010011101111101010011001001010001100111010010000010100010101001010111100101001010000000001000101110100100101110010010111101001001;
		5'd25: 256'b1100000110110101001011111010011000001011101110001010110101010110100010111001110011010100001011001100010101110100010010101000000111101010000101011010000110011110000000010011000101010001111011000110000011111001101111000101111000011010001011001110011101101110;
		5'd26: 256'b0000110111011011000111010100001110011101011000011000010111100111111011111111100101101111100100001101100100000000101001111000010000001111011000011111100000000111111111111000111001110011100110100110111010111110100100101011101111010110110011000001110011100010;
		5'd27: 256'b1100001110101011100111101110101010000000111111100011110011011111011001000100010101111010000011001010111010011110110110111101010011001000111001100000110010000011110000000001100101110101011000001001111111110001111000110110011111000111111111111111010000111100;
		5'd28: 256'b1100000011000001111100011110010011101110000110110010110110000100001110100101111100101111000000000000011101100110101010010101001110000011001000111100101101100101100001100111111110001000000111010111110110000111100110100101000111011101101100001011100100010011;
		5'd29: 256'b1111111010110111110001100000100010000011110001001100111011010111110110100011000011110011001101110011011000010001101110111001011110011011001101001111101101101101011001101001100001000001101100000001011010111101001101111000111000000101000010000010011110111011;
		5'd30: 256'b1110001110011011100010001000000111100111010111100010110010100001111110111111111001101110001111010111010000111010110101111100010111001110010010011001000000011111100011001011001011101100000101100101011110100101111111010011111001010011111110111000100111111110;
		5'd31: 256'b1110100111110010010101100101101100101011010010111101100001001100010000111100100010101111111110001100110100110100110110010100010000010101000011101001010100101001001101101011001001001110011011101101110101101001110100001111001011000001101111011001010111111000;
	endcase;
	return out;
endfunction
function Bit#(64) get_prev_enc_page1(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b0000110010000000000000000000000000010100100100000000100001000000;
		8'd1: 64'b0010000000000000000000000000000000111000010000100000100001000000;
		8'd2: 64'b0000000000000000010000000110000000000000011000000010100000000000;
		8'd3: 64'b0000001000000010000001000000000000001000100010000010000100100000;
		8'd4: 64'b0101000000000000000001010000000010000000000000000000000011000000;
		8'd5: 64'b0000001000110000000000001100011000000000101000100000000000100001;
		8'd6: 64'b0001010010010100000000000000000000000000000000000000000000000000;
		8'd7: 64'b0000000000000100000001000001000000000000000010000100000101000000;
		8'd8: 64'b0100000000100011000000100000000000000100000100000001001000000000;
		8'd9: 64'b0100011000000000000000001000000000000000000000101000000000000000;
		8'd10: 64'b0011000100010000101000001001000000000100000000000000000000001000;
		8'd11: 64'b1000000001000001000000000000000000000000000000000010100000000001;
		8'd12: 64'b0000010000000000000000000000000000000001000100000010000000000010;
		8'd13: 64'b0000000000000000000000000000101000000001110000010010000000000010;
		8'd14: 64'b0100100000000000100000000000000010000000000000110000001000000101;
		8'd15: 64'b0010000000000001000101000000000010000000000000000010000010000000;
		8'd16: 64'b0000000011000000000000000000000011100000101100000000000000000001;
		8'd17: 64'b0000100000000000000000000001000100001000000001000001000001000000;
		8'd18: 64'b1000000010000000001000100000000000000000000000000000011000100000;
		8'd19: 64'b0100101000010001000010100000000010001000100000000000000000000000;
		8'd20: 64'b0000000000000000000000100000100100000000000000010000001001010010;
		8'd21: 64'b0000000111000000100000000011000100000011000000000000100000100101;
		8'd22: 64'b0000000000000000000001000000100000001000000010000000000000000000;
		8'd23: 64'b0000110000000000000000000000000000010000000000010000000000100000;
		8'd24: 64'b1000000000110010100000000000000000000100000000000000000110000001;
		8'd25: 64'b1000001000000000010000100000000100001010000000000000000000000000;
		8'd26: 64'b0000000010000101000000010000000000000011000000010000010000000001;
		8'd27: 64'b0000010010000100000000010000000000000000000000100000000100000010;
		8'd28: 64'b0000000000000010000100000000000100000001000000000000001000000000;
		8'd29: 64'b0110000010000000000100000000000000000000010000000001000000000000;
		8'd30: 64'b0000000000000000000000100000000000000000000001010000000000100000;
		8'd31: 64'b0000000100000010000000001110000000001000000001100000000000000000;
		8'd32: 64'b0000000001010000011000000000100000000000000100000000000000000000;
		8'd33: 64'b0000000000010101001000000000001000000000010000001100000000000000;
		8'd34: 64'b0000000100100000010000000100000100010000000101000000000000100001;
		8'd35: 64'b0000000100010000000000000000100000000000000000001000001010000000;
		8'd36: 64'b0000001000000000100101010000001000001000010000000000001000000000;
		8'd37: 64'b0110000010000001000000000000000000000000110000000001000000000100;
		8'd38: 64'b1000000001000000000000000000001000000000000001000000000000010100;
		8'd39: 64'b0000000010000000000010000001000000000000100000001100000000000000;
		8'd40: 64'b0100000000000000000000000001000000100000010001010000010001000000;
		8'd41: 64'b0000000100010000000000110000000000000000000010000001000000000000;
		8'd42: 64'b0000000000000000000000000000100000000000000000000100000000100000;
		8'd43: 64'b1001000110000000000000000000010000000000000000000001000001000000;
		8'd44: 64'b0101010000000001001100100000100000000010100100010000000000010000;
		8'd45: 64'b0000100000000000110000001000000000000010000000000000000010010010;
		8'd46: 64'b0000000000000000000000000000000100000100000000000100001111000000;
		8'd47: 64'b0100100000000000000010000000000000000000001000000000000010010000;
		8'd48: 64'b0000000000100000000000010000000001110000000000001000000001001000;
		8'd49: 64'b1000000000000001001000000000000000000000100100010000011000000000;
		8'd50: 64'b0000000000001111000000000000010100001000000001000000000000000000;
		8'd51: 64'b1000111000000010000010000000000000000000000000001010000000000000;
		8'd52: 64'b0100010000000000000000000000000000000010000001001000000000010000;
		8'd53: 64'b0100000000010100010000010000000000000000000000000000000000000000;
		8'd54: 64'b0100000000000000000000010000000000100000100001001000000001100000;
		8'd55: 64'b0000000000000010110000001100000000000000000000000000010000000000;
		8'd56: 64'b0000000100000001000000000000000001010000000000000101010000000001;
		8'd57: 64'b0100001000000000000000010010000100000010000000010100010001000000;
		8'd58: 64'b1000000001000000000000000000000000000010000001010010001000001101;
		8'd59: 64'b0000000000101000000010100000000000000000000000000001000101000000;
		8'd60: 64'b0000000100000000001000001010000011000000000000000010000000000000;
		8'd61: 64'b0000100000000000000100000101000000001010111000000101101000100000;
		8'd62: 64'b0000010000000010000000001000000001000010000000000100001000000000;
		8'd63: 64'b0000000000010000001000000010000000001000000000000001000000000000;
		8'd64: 64'b0100000101000000100010000001000000001000100000001000010000000000;
		8'd65: 64'b0000000100011000000000001001000000000000000100000000000000000000;
		8'd66: 64'b0000000000000010000000000000000000010000000000000011000100000000;
		8'd67: 64'b0000000100010000000001100000000000000100000000001010000010000100;
		8'd68: 64'b0000000001000000010000100010000000000000000100000000000001001000;
		8'd69: 64'b1000010000000100000000000000000000000100000101100000000000000000;
		8'd70: 64'b0000000000000000000101000000000000010000010000000100100000001000;
		8'd71: 64'b0010000110000100010110000000001000010010000000000000001000000100;
		8'd72: 64'b1000000000000111010000000000010000000000000100000000000000000000;
		8'd73: 64'b0000000000000000000001000000111000000100000000000000000011000000;
		8'd74: 64'b0011100000000000000000100000000100000010000000001000000000000000;
		8'd75: 64'b0001000010000000000000010000000000000000100001001000000000011000;
		8'd76: 64'b0000000000000000000000010001000100000101000010110001000000000000;
		8'd77: 64'b0000000000000000100010000100000000010000000100000000001000001000;
		8'd78: 64'b0000000000001010000000010100010100000000000010100110000000000000;
		8'd79: 64'b0000000000000100000000001000100001100000000011000000000000000000;
		8'd80: 64'b0000010000000000000000010000010001001000000100011000000001000100;
		8'd81: 64'b0001000010000000000000000000001000011000000000000000000000000000;
		8'd82: 64'b0000000000000000001000000000001000001000000000100000100000100000;
		8'd83: 64'b0000000000000001100001000100000100100000000000010000000100000000;
		8'd84: 64'b0000001000001000100000000100000000000000000000010001011000001000;
		8'd85: 64'b0000001000010001000000000000000000000100100001000000000000000000;
		8'd86: 64'b0010000101000000000011010000000010000010010000000000000100000000;
		8'd87: 64'b0001000010010000000000000000000000000000000010000000010000100100;
		8'd88: 64'b0000001010000010000010010000011000000000000000000000010100000000;
		8'd89: 64'b0001000000000000001000000000001000000000000000000000000100001000;
		8'd90: 64'b0100000000000100000010000000000010110000000000100000001000000000;
		8'd91: 64'b0000000000000000000000000000010000010000000000000001000000000001;
		8'd92: 64'b0000100000100000000000000000100000000010110010100010000000010010;
		8'd93: 64'b0000000100000011010000000001100000000000000100000000000000100010;
		8'd94: 64'b0000000000000000000010000000000000100000000000000000001100000000;
		8'd95: 64'b1000000000100000001100000000010000100000000000000000000000000000;
		8'd96: 64'b0000000010000000000000010010000000000000000000000000000000000000;
		8'd97: 64'b0000000000001000001000001000000000000000001010000010000000000001;
		8'd98: 64'b0000000000000000100000100001000100100000000000100100010000000000;
		8'd99: 64'b0000000010000100000000000100000100000000000000001010010000000000;
		8'd100: 64'b0000100000000001100000011000100100000000000000000000000010100000;
		8'd101: 64'b0011000100100000000000000010000001010000000001000100000000000000;
		8'd102: 64'b0000000000000100010000100000010000001000000000001000100000000010;
		8'd103: 64'b0001010000000000000000000010000000000010001000100100001000000010;
		8'd104: 64'b0000001000000000000100000000000000010000010000011111000001001001;
		8'd105: 64'b0010000000000000000000000000001000000000000000010000000000000000;
		8'd106: 64'b0000010000110000000000000001000000000100001100010000000010000001;
		8'd107: 64'b0000000010100001000001000001000010000001000000000000000000000000;
		8'd108: 64'b1000010000000000000100100000001000000000000000000000100100001000;
		8'd109: 64'b0000000010000100000010000000000000000000001000010000001100000011;
		8'd110: 64'b0000001000000010010000000000000001100000000110010001000000100000;
		8'd111: 64'b0001000000000000000000010000000001101000000010001000000000000000;
		8'd112: 64'b0101000000000000000100000001000000000000000001001000001000000000;
		8'd113: 64'b1001000000001000000000001000000000000010000001000000000100000000;
		8'd114: 64'b0100001000000000001100000010000000000000000000001001000000000010;
		8'd115: 64'b0010100000000000000001010000100100000001000000000000000000001011;
		8'd116: 64'b0000000000001000001101000001000110001000000000000001000100000000;
		8'd117: 64'b0000000100000011001000000010010100000100011001000000000001000010;
		8'd118: 64'b1010000000000000000001000100000000000000000000000010000000000000;
		8'd119: 64'b0000011000100000000000010000001100000001001001001000000000000000;
		8'd120: 64'b0010000010010001010101000000000011000000000000000000010000000000;
		8'd121: 64'b0000000001010000001010000000000101001000000000000000100100010000;
		8'd122: 64'b0000000000000000000000000000000000000000001110010001000000000000;
		8'd123: 64'b0000001000000000000000000000000000000000000000100000000000000000;
		8'd124: 64'b1000000001000000001000000001000000000100000001100000001010001001;
		8'd125: 64'b0000000000010010000000000000010010000000000000000000000000100000;
		8'd126: 64'b0000000000000001000000010000000000010010000001100000010000000000;
		8'd127: 64'b0100000000000000000000000000000000000000001100010000000000100000;
		8'd128: 64'b0000000000110000000111000000000001100100100000001100000100100101;
		8'd129: 64'b0000000110000000001000001000010100000000000001000010000001000000;
		8'd130: 64'b0000000000000001000010000000100000000001000001000001000000100000;
		8'd131: 64'b1000000000100000000000000000000010000000000000100100000000000000;
		8'd132: 64'b0000000010000000000000000110000010000000000000010000000000000010;
		8'd133: 64'b0100000010000000000000000000110000001000000000000000000000000100;
		8'd134: 64'b0011000000101001000001010000000000010000000000100000000001000100;
		8'd135: 64'b0100000000000000000000000100000000000000001000001000010010010000;
		8'd136: 64'b0000000100010000000000010000110010001000000000000000000000010100;
		8'd137: 64'b0000100100100010000000001001000000010000100010000000100000010000;
		8'd138: 64'b0010001100000100000000000100000000000001000000100000000000000000;
		8'd139: 64'b1000000000000100000001001000000010000001000000000010000101000000;
		8'd140: 64'b0011000000000000100100000000000000000000000000001000000000100000;
		8'd141: 64'b0001010010000000010000100010010010000000010000000000000010000000;
		8'd142: 64'b0000010010001000000000010010100000000000000000000000000000100000;
		8'd143: 64'b0000100000000000000000000010000110000010000000000000000000010100;
		8'd144: 64'b0000000010000000010000000000000010100001000000000000000000000100;
		8'd145: 64'b0000000000000000010001100000000100010001001000000000000000010000;
		8'd146: 64'b0000001000100000000001000000000000000000000000000010000000000000;
		8'd147: 64'b0000000000000000010000000010000001000010100000000000000000000101;
		8'd148: 64'b0000001001000010000000100000000000000001001010000000000000000000;
		8'd149: 64'b0000000000001000000000000100000010100000010010100000000001000000;
		8'd150: 64'b0010100000000100001000010010000010001011000000000000011000000000;
		8'd151: 64'b0010000000000100100000000000100100000000000000101100000000000000;
		8'd152: 64'b1010000000110001000000010000000000000000001000000000000000000000;
		8'd153: 64'b0000001000000000010000000010000000000000100000100000000100000010;
		8'd154: 64'b0000000000000000000101010100000000000010100000000001001000000000;
		8'd155: 64'b0000000010110000000000010000010000010001000000000001001100010000;
		8'd156: 64'b0000000000010000000000000000100000000000100000000000000000000100;
		8'd157: 64'b0010000100000000000000000000000000000000000000000000010010000100;
		8'd158: 64'b0000100000000010000000000000000000100000000101000000001000001010;
		8'd159: 64'b0010000010000110000100000000000010010000101100001000011000001000;
		8'd160: 64'b0000000000000000000000000011000000100000000000000010000000100010;
		8'd161: 64'b0000000000100000000000000000100000000000001000000000000000010000;
		8'd162: 64'b0000000010000000000000000000000000010000100000110000000010000010;
		8'd163: 64'b0000000100000100000000000000100000000000000000000000000100000000;
		8'd164: 64'b0000000000000000000000000000010000000100001001000000000110111100;
		8'd165: 64'b0000000000000000010100010000010100000000101000100000000000010000;
		8'd166: 64'b0000000000000100001000000000000010100001100000010001000000010010;
		8'd167: 64'b1000100000000000000000000000001011000000000000010010010001000000;
		8'd168: 64'b0000000000000001000000100010000000000000000000000000100101000000;
		8'd169: 64'b0010010010100000000000000000000000000000011000000100000000000000;
		8'd170: 64'b0000100000000000000000000011010110000010011000001000110010001000;
		8'd171: 64'b0010000000001000000000000010001100000100100000110001000001001000;
		8'd172: 64'b0000001000000000000000000000100000000000000000000000000000000000;
		8'd173: 64'b0000000000000100011000000000010000000000011000000000001000000000;
		8'd174: 64'b0001000000000000000010100000000100000001101000000001000000010000;
		8'd175: 64'b0100000000010000000000101000000000000000000000000001000000000000;
		8'd176: 64'b0000000000000100000010000000000000000000000000000010010000100001;
		8'd177: 64'b0000000000010100000000100000000010000000000000000000000001001000;
		8'd178: 64'b0100010000100000000100000000000000001000001010100000000000010001;
		8'd179: 64'b0000000100000010000100001000100100000000100010000000000000000000;
		8'd180: 64'b0000000010000000100100010000000000001010000000000000001000010000;
		8'd181: 64'b0010000001000000000000000000000000100000010000000100000000010000;
		8'd182: 64'b0100000100000001000000000000000000000010000010000010000000000001;
		8'd183: 64'b0000001001000000000000010000001000000000101000001000000101001000;
		8'd184: 64'b0000000001001001000010001011100001000000000001000000001000000000;
		8'd185: 64'b0000001101000000010100000001010000000100000000000000001000000000;
		8'd186: 64'b0000000000000010000001000100100000000000000000000000010000000000;
		8'd187: 64'b0000011100000000110100010000000000000000010000000000000000100000;
		8'd188: 64'b1001000000001000100000000001000000000000000000100010100100000101;
		8'd189: 64'b1010000000000000000000000000000000000000010000000000001010000100;
		8'd190: 64'b0000000000000001000000000001000000000001000010000000000000000000;
		8'd191: 64'b0001000000000000001000000100000000100000010000000000100101000000;
		8'd192: 64'b0000000000000000000000010110000010000000010000000000000001000000;
		8'd193: 64'b1100000001001000001000000000000000000100000000010000001000010000;
		8'd194: 64'b0100000000000000000101010000000000000000100001000000000000100000;
		8'd195: 64'b0100001110100000010000000000001011000010001000000000000000000000;
		8'd196: 64'b0000011000000000000101000000000000001000000000000010000100010100;
		8'd197: 64'b0010000000001101000000100001000001000000010000000001100100001000;
		8'd198: 64'b0000000000000000000001100001000000000000000010010000000000000000;
		8'd199: 64'b0000000001000001000000000000000010000000100000000100000010001000;
		8'd200: 64'b0001010000100100000000000000110100001000000100000000000000001000;
		8'd201: 64'b0000001100100000000000000000010000110000000001000000001000001000;
		8'd202: 64'b0000000000000100100000011000010000000000000000100000000000000000;
		8'd203: 64'b0000000000100000010000010000000000001000000000010000000001000000;
		8'd204: 64'b0000000100000000000001000010000000100001000000100010000000100010;
		8'd205: 64'b0001000000000000000000000000000010100000000000000000000100000100;
		8'd206: 64'b1000000000000000001001000000100000000000000000000000100000000010;
		8'd207: 64'b0010000000000001000100000010011010000000000100000001000101000011;
		8'd208: 64'b0100000000000000010000100000000000000000000000000100000000000000;
		8'd209: 64'b0000100000000100000000010000100000000000000010001010100010000000;
		8'd210: 64'b0000000000000000000010000000000101100000001000000000010000100000;
		8'd211: 64'b0010000000000000000000010100000000010000000000000010100000000100;
		8'd212: 64'b0000010100000000000000000010000001010100000000000000000001000000;
		8'd213: 64'b0001000000000000001000000000000000100010000000001000100001010000;
		8'd214: 64'b0001000010000000100000000000000000000110000000001000001000001000;
		8'd215: 64'b1000001001000000000000100000000000000000100000101000000110000000;
		8'd216: 64'b0000000000000000100001000000000000000010000000010001000000000000;
		8'd217: 64'b0101000001000000000000000000000000000000000000000001000000000001;
		8'd218: 64'b0010001000011000000000001010000000000000100000000000100001010000;
		8'd219: 64'b0010000000000000000000010000000000100000000100000100000000000000;
		8'd220: 64'b0000000000000000001000001000010000010000010000000000000100000100;
		8'd221: 64'b0000000010000000000100000000000010010010001000000000000000000000;
		8'd222: 64'b0000001000000000001100000000000100100000000000000000000000010110;
		8'd223: 64'b0000000010000100000000010000000000000001000100000100000000000000;
		8'd224: 64'b1000001000010000000000000010001011000000110000010000110000000010;
		8'd225: 64'b0000000000001000100000000000010010000100000000000001000000100000;
		8'd226: 64'b0000000000000000000000000000000001100001010000000001000010000000;
		8'd227: 64'b0000000000100000000000000000000000000100000000000000100000000001;
		8'd228: 64'b0000000000000000010000000101100000000100010001001000000000011100;
		8'd229: 64'b0000000000010000000010000001000000000000000000000001000100000000;
		8'd230: 64'b0000000000000100000000000000100000000001000000001010001001000000;
		8'd231: 64'b0000011000000000000001010000000000000000000000010000000000000000;
		8'd232: 64'b0000001010000000100000000000000000000000000000100000000000000100;
		8'd233: 64'b0010000000000010000000000000000000010101000000000100000000011100;
		8'd234: 64'b0000001000000001000000000010000000100100000000110000000100000000;
		8'd235: 64'b0100000100000000000100000000001000000000000000000000001010000000;
		8'd236: 64'b0000000000000000000100000000100000100000000000000000000100000000;
		8'd237: 64'b1000000000000000000000000000001000001000010001100000000000000000;
		8'd238: 64'b0100010000000000001000000001000000100111000010000000000000001000;
		8'd239: 64'b0000000010110000000100000000000100000000000000000000000000001001;
		8'd240: 64'b0000001000000000000000000101000100000000101000000000000000101001;
		8'd241: 64'b0000000000000000000000000000001000001000110001000000000000000000;
		8'd242: 64'b0000000000010000010001101000010100100000000010000000000000000001;
		8'd243: 64'b1010000000000100000010000001100001101000000000000000000000000000;
		8'd244: 64'b0100000000000110000000000000010000100000100000000000000000000000;
		8'd245: 64'b0010000000000000000000000000001000010000000000010001100000001000;
		8'd246: 64'b0000000000000100010000000000000000000000000000010000100000100000;
		8'd247: 64'b0000000000000000000100010000000000000000000000000000000000000001;
		8'd248: 64'b0000000001100100010000000000001000000000000000010000000000000001;
		8'd249: 64'b1110000011000110000000000010000000000000000000000000000000001000;
		8'd250: 64'b0100100000100000010001000000010000000000000000001000000000000000;
		8'd251: 64'b0101000000000000000000000101001000000000100100000010000000010100;
		8'd252: 64'b0010001000000000001000000000000000000000000000000001000000000000;
		8'd253: 64'b0000000000000001000000000000100000000000000000000000000010000000;
		8'd254: 64'b0000100001010000010000000010000010000000100000000001000001000000;
		8'd255: 64'b0000000000000001000100000000000000000000000000010000000101000100;
	endcase;
	return out;
endfunction
function Bit#(256) get_msg_bit_page2(UInt#(5) counter);
	Bit#(256) out = case(counter)
		5'd0: 256'b0011100010000001110110011011110100111110001110001011001110001111100110010010111110001101101101001100010001101011100010101101000000110111101001000001100111111001010001000110010111010111111111100011001111011010101101101000100001010010000011110110001000011111;
		5'd1: 256'b1001010000100110001100110100010110010000111100101111010100000000111011100010000111110100001000000100010001110011111100110100010110010000010010010010000101100111000010010010111001101010111011000000010101010101110011011111110010111111011111111011101000000011;
		5'd2: 256'b1100011110101001111010011011101000100101100100001001111001110011000111001001001000101100111101101010101010110010111010100110100010110110111010000001010010111011111110001010011110101111110001111000011001001111010011111010001010100110111010100010100011010001;
		5'd3: 256'b0101011110100111101111110011001111100110111100100010111011000100011011110100011000001100010100101011011000111111111000000100000100100010100011100111001101101000101000101011111111000001000101101011100010001111101011011010100000111010111011101011101111110111;
		5'd4: 256'b1000000011010011101100001000101011110100000000010000101000101110011101101010001000011000111110101000001011010001110101110110100010001110001101110011001101110010010001001110111000010100011110011001010100010111111010001101100111111111101100000110011011110011;
		5'd5: 256'b0111101101110101000100001110101110001100100110000110001011110111110110000001111011110011110011000011001100010110011101010110100000100111001010010111001010010111010001010100001101101111010101100100101100001101000111111111101111101000110010111111010100001000;
		5'd6: 256'b0011010001100101001101110000100111110011101000001101110110110000101100001000111010101011100100001010100001101010111001001011111000010011000111111100010100101001000100100011111101011100101110000011111001101001101001000001011011100000010001000011100000010101;
		5'd7: 256'b1100101111001011000101100100010100001110110111000011011101011101101011100001011111101010111110110101100100000101010010111000101111111001100111011010100101100011001000001011000110101101111111010110001011110101100111100001110110000011101011000010101010110110;
		5'd8: 256'b0000001000101100110000000110010000111001010010000111000010000010010101001011110000100100001101001011001011011110011001111100111111101001111010111111111011111100111101001010110101111101100011111000011001111001001000000000110010010100010101001000001001101011;
		5'd9: 256'b1100100111010101110100010000011101000001000000010001001011100001001101011110011110001010010110100001101101100010100010111110011101010101111111110100011010110000111111100000111010111111110000000110011111001100110100111111000010001010110100110001101111010110;
		5'd10: 256'b1101000000011000100000100010011001010000110101100101100011001001001101110110100111010110110100010101000101110110011101111101101101000100100110011110011000001010110000001011001011100010010011110001101001010110001110011100000111100110001110110111101011111111;
		5'd11: 256'b1010010001111101110110100100100001010101101000011111101100110001111011100011011010011001001001101010010100001000101000101110101011000100011000011101011111001001101011000011011111111010101011011001010010101110110011001100100110111101000010011001101011011101;
		5'd12: 256'b1110101100101101001001111101100010000011100001011001001110100000111011000100100101111010000110000110101010110101001010011000001000110101110011101100110010101101110101001011000110110001010011001001110000100110010001001101110100001100101000101111100000010000;
		5'd13: 256'b0100100100100111110111001100101101110101001100101010000111111111101110100001011100011011010011110001011001100010011000110011011010000011011110111011001101101111110001100000110000111001000111110000111001011001011110010111000110011111100010000110011011000000;
		5'd14: 256'b0011000000001000001111100001001111101011001011111010110011101010111111000100101111110010011110001010110011111000100101110011111101001010101001001011101000000100010011010110101000100100101001010110010111111010000011111110010111100100111110110101000100000010;
		5'd15: 256'b1110010000110101101101010001010011010011110011110011101000010000000111110101100001101110110101001100011111111010011101011110011101000111000111010001010100000100111111011100111001100100011001000110101000001011000110001111110010110000010000010000110100010111;
		5'd16: 256'b0101010110010110010010011010001100010101010001001000111010001010011011011101100110100101100100010001110001101011001010100000001010110001001111011101110100101010010111010010010100001001110000101010000111011111100100000001101000110001110111110000110110111011;
		5'd17: 256'b1001111001101010111010100110010000100111111111011101110100110111001010110110001010110110101000110110010010110110011111111000011000010011010110001110101000001010010000111111001011000010100100101111110001101010000010011101011101001010010100000000110000110001;
		5'd18: 256'b1100011001001111010000110110111100110110101100100101110100011000101101000110001100011000101100110111000000100000011111000111011010001110001110010010001111100111011010001001000001000111101011010111101011001011010000011000111000101111110011000110011000110000;
		5'd19: 256'b1011100001100101111000100000100111110011000111111100001110110010001010101101110000101110010000101110011011110111011010111111100000110001111111110111001111001011010101110000000011100101011001001010001101110010100111001111101111001111110010001011000101101101;
		5'd20: 256'b1111110011010001101100010100010000000101111011010100000000110100111111001001000100010010000011001010011011010000011100001110010101010101000001001000100100000110101110111000001100011101010001000001111001011001100100111100111100001001000010001011111010100011;
		5'd21: 256'b1100101001011010100110010010000110111101011011111100101110001011010011010010100101110011110111001110101101010111111001001110011100100011011110000100000100111110110100101100001010110101000100001001110100010100110110010010100001010111101101110001110110001101;
		5'd22: 256'b1101000000011110111101000001101111110000001110100110001111000001000111001110111101101001011100001001000110111001001100010001000011000110111011101110010111111010000101110110101100010000000111010111110111010001000011001011101101011100111000101000110001000111;
		5'd23: 256'b1010110111010000110101101111110011110110011110010110011000011001001000001111101011111000101101110010111100010001111100111000101011100000000101010110110101100110100001000110100101101011111110010101001111000110000111001010111111110001101011011000011111001101;
		5'd24: 256'b1101110000100111111011000011000110001100011000000000000101010110100011000101011000000111100001001011000010110110010110101001110000011110000000011011011011000111111100011100000001101111000000011010110010111101110110110011101001100000110100000011011101000010;
		5'd25: 256'b1100111100101111110010100110111111010000111101101111101100000000001011010000110111001000011010010110111111110100011101000010011010111111111011000100000011100000001101110111110011000011001111111111000011010000100100100111001000101100010000100101000001110100;
		5'd26: 256'b1101000011100111110110100110011000111011110011100001001110111101000100000010101001100110001110000100111001100010100100011111101111110110001101111100101000000010110101000000101111101111100000101110000010100111000101110111001001110011001000110010111111001000;
		5'd27: 256'b1110010011010111010111101001101110001101010010110001000000110010101001101110100011011110000001000111110110011111000101111010000101001000101110000000010001100010100100010110110111000001101111000101100111001111111011000010001101011111010010011011000100010010;
		5'd28: 256'b0100111111111101101101101110111100010010101101011100010101110101111000111010100000101101110000111101011100010100110011001001111110111111010100111011110000000000010111010110110111110100011011100001011100011010100100101000111100110011100110010101101010110010;
		5'd29: 256'b1110101111111010100010011101100111011010101000110101100011110111000000000001110110111001111100100010000001100001110001001011111000100111101100101010001010001011110010001010100101010000010111101111010101000000011011111110100110010100001010101001101000010001;
		5'd30: 256'b0000111101001100101010011111111010001101001011110100011001101011000011010011010011010111110011000111100010101000111001100111111101110010001011000111111100001110101000001000110010111110101100001101010111010011110100100101110000001101001011110010001110011001;
		5'd31: 256'b1111010001100101000011101100011010010001100010100001110011110100011011010100000111100100001010011101100001011101111110011101000000110100011110101011011100100110110101111110000110010011111100101000101010011000001110111110010101001000010010001101110011101101;
	endcase;
	return out;
endfunction
function Bit#(64) get_prev_enc_page2(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1000110010001011010000001000000000011100100100100001100001000000;
		8'd1: 64'b0010001010011000001010000000000000111000010100100000100011000000;
		8'd2: 64'b0000000000000000010000000111000001000000011100010010101000011101;
		8'd3: 64'b0001011010110010000001100001000000011001100011000010000100111001;
		8'd4: 64'b0101000000000001000011010000000011000000000000000000001011000000;
		8'd5: 64'b0000001000111000000010001100011000000000101100100000010000100001;
		8'd6: 64'b0001010011010100001001001100000000101000000000000000000001010001;
		8'd7: 64'b0000000111010100000001100001000000010000000010000100100111010000;
		8'd8: 64'b0101010000100011000000110010000100000100010100000001101000000010;
		8'd9: 64'b0100011000000000001000001000000100000000000000111000100010000000;
		8'd10: 64'b0111000100010000101001001101011010010100000010000000100000001000;
		8'd11: 64'b1001000001000001000000000010000000010001010100110010100000001011;
		8'd12: 64'b1010010001010001000000000000100000000011000100000010000000000010;
		8'd13: 64'b0000010000000010001000000000101000001011110010010011100000011010;
		8'd14: 64'b0100100000010010100010000100000011010000000000110000001000000101;
		8'd15: 64'b0110110000000001000101000000000110010000100000100010000010000000;
		8'd16: 64'b0010000011001100000000010001001011100000101111000100100000000001;
		8'd17: 64'b1010101000000000000000000101000100101000000001000011000001000000;
		8'd18: 64'b1000000110000000001111100000000000110000000000001000011000101000;
		8'd19: 64'b0100101000110011000010110100000010011010110100011000100000000000;
		8'd20: 64'b0010000000001001001000100000101100000001000001111000001001011010;
		8'd21: 64'b0011000111110000100010001011001110000111010000111000100010100101;
		8'd22: 64'b0000000001110010000001100000110001001000001010000000000001000001;
		8'd23: 64'b0011110000011000100000100000000000110101100010010010000100110000;
		8'd24: 64'b1000010100110010100100000011100000000101101001001000000110010011;
		8'd25: 64'b1010101010000001010000100101001110001111001100100010000000100000;
		8'd26: 64'b0001001010010101000001010000100001001011110000011000010000001001;
		8'd27: 64'b0000010110000100000000010000000000100000100000100100000100000010;
		8'd28: 64'b0100100000000010000100100000011100000001010010000000001010000010;
		8'd29: 64'b0110000010100001000100000000000010000000010000010111000010000000;
		8'd30: 64'b0100010010000001000000100000001000000000000001010000100000100000;
		8'd31: 64'b0000000100000010100000001110000000011000100001100100001011000000;
		8'd32: 64'b0100000001010000111000001001100000010000001100000000000000001000;
		8'd33: 64'b0001000000010101011001000010011000000000010100001110000000100000;
		8'd34: 64'b1001000100101000010000010100010100011000000101001000000001100111;
		8'd35: 64'b0000101110010010000001001000100100010000100000001000001010010001;
		8'd36: 64'b1100001001000000100101010100001100001001010000000100001000100001;
		8'd37: 64'b0110010110000001000101010000000000100011110000000001000010000101;
		8'd38: 64'b1000000001000101100100000001011000000100010011000010000000010100;
		8'd39: 64'b0000101010001000100010100001000000000010100010001100000000000000;
		8'd40: 64'b0110000100000100000001000011100010100000010001010000010001000000;
		8'd41: 64'b0000000101010100000000110010000000000100000010001001000000000010;
		8'd42: 64'b1000100100011000010000000000100000000010000000000110000100100000;
		8'd43: 64'b1001100110000100010010000100010010010000000001000101000101001100;
		8'd44: 64'b0101011000010101101101100001110001000110110100010001000000010000;
		8'd45: 64'b0000100010000001110000001001101100000010001100010100000010010010;
		8'd46: 64'b0000000000000000000000000000000100000100001000010100001111000000;
		8'd47: 64'b0100100100011101001010000000000000000000001001000010100010110000;
		8'd48: 64'b0011000000100000000100010001010001110000000000011000000001011001;
		8'd49: 64'b1000001100000001111010000000000000000010100100010000011000010100;
		8'd50: 64'b0000000010001111000000000100111100001101000101000011000100010000;
		8'd51: 64'b1010111010000011000011010000000000100100111000101010010000000000;
		8'd52: 64'b0111010000001000000100010010000000000010000001011000010000010000;
		8'd53: 64'b0100000000010100010000010000000000000000000000000011000000110000;
		8'd54: 64'b0100000000100000000000010101000000110001110001011010010001110001;
		8'd55: 64'b0000010001000110110000001100001000000000000000101100010000010000;
		8'd56: 64'b0000001100000001011001000000000001010000000010000101010011000001;
		8'd57: 64'b0100001000001000000001010110001100000010000011010100010001000100;
		8'd58: 64'b1000000001000011000000110000000000000010000101010010101000001101;
		8'd59: 64'b1000000000111000000110100000001000001000000010010011001101000011;
		8'd60: 64'b0001010100000000001001101010010111000011000000000010000010100100;
		8'd61: 64'b0000100000100001010100000101000011011110111000000101111100100100;
		8'd62: 64'b0010010010000110000001101000000001100010000001001111001000000000;
		8'd63: 64'b0000110000010000001001001011000000001100001000000001010000000000;
		8'd64: 64'b0100000101000001100010000001000100001100110000011000010000010011;
		8'd65: 64'b0000000101011000000010001101100110110000010100001000000010000000;
		8'd66: 64'b0001010000000010000000000000000000010000000000000011000100001000;
		8'd67: 64'b0000001100010000000101100001000001000100000100001010100010000110;
		8'd68: 64'b0000100001100010010000101011110001100000000100100100001001011000;
		8'd69: 64'b1000010000100100000000000010000000100110001101100010100000010010;
		8'd70: 64'b0000000000000000101101000010000000010000010101010100100000001000;
		8'd71: 64'b0011000110000100010110000000001010010011000000100001001100010100;
		8'd72: 64'b1010000100100111011000000001011010000000000100001000001000000010;
		8'd73: 64'b0000100000000000000001000100111000010100000000000000010011000000;
		8'd74: 64'b0111100000100000000000101000000100001110000000011101000001000001;
		8'd75: 64'b0001010010011100000000111100100001000000100001001000000000011000;
		8'd76: 64'b1000010000000010100101010001010100000101000110110001011000000000;
		8'd77: 64'b0100000100000000100010000100000100010000000101010000001110101000;
		8'd78: 64'b0010011010101110000001010100011100000000000010100110100000000010;
		8'd79: 64'b0101100000001110000010111000101001100000000011000000011000111001;
		8'd80: 64'b0100010000000101000001010010010001011000000100011000011101001100;
		8'd81: 64'b0001100010100000000000000000101010111100000001100000000010000001;
		8'd82: 64'b0100000000000000001000000000001000001100000000110111101000100000;
		8'd83: 64'b0000000100000101100101000100010101100011100000010001100100000000;
		8'd84: 64'b0000001010001000100000101110010010000000100000010001111001101000;
		8'd85: 64'b0000011000010001000000000000000000000100110001000000010000000000;
		8'd86: 64'b0010001101000000000011110000011010000010010101000000000101010101;
		8'd87: 64'b0001000011010010100000000001000000000001000110000000010000110101;
		8'd88: 64'b1000101010000010000010010000011100000000001000110000010100000000;
		8'd89: 64'b0001000000100100001000010010011010100010000000010100000100001010;
		8'd90: 64'b1100000001000110000010000000010011110000000010100001001000001001;
		8'd91: 64'b0001000000000010000110000010010000011001000000000001000010000001;
		8'd92: 64'b0000100100101010000000001001100000001011110010100010101010010010;
		8'd93: 64'b0000000110010011011010000001100000101000010100010000100011100010;
		8'd94: 64'b0010100000000001000010000011000001100000000001000000101100000000;
		8'd95: 64'b1000000100110001001100000000010000100000000000000100000000000000;
		8'd96: 64'b0000000110100000010110110010101000000000000001010010010011101100;
		8'd97: 64'b0001000100101000001100101011000000000001001010100010100000000001;
		8'd98: 64'b0010000000000010101000100001001101110010000000100100010000000010;
		8'd99: 64'b0000000110000110001000000100000110010000001000001010010000000000;
		8'd100: 64'b1001100100001001100100011000100101011101000000001001000010100100;
		8'd101: 64'b0011100100100000010000001110010101010000000001100100000100000100;
		8'd102: 64'b0100000000010100011110100000011001101000101001001000100000000010;
		8'd103: 64'b0001010001000000000010001010000000000011001000100100001000000010;
		8'd104: 64'b0000111000000000000100000000000000010010010000011111110001001001;
		8'd105: 64'b0010001000000011001100000000001000000000000000110010010000000000;
		8'd106: 64'b0000111000110000000010000001000000100100001100010000000011010001;
		8'd107: 64'b0000000010100001000001100001100010010001000000000000000000000000;
		8'd108: 64'b1000011100000000000100100000001000010001000011001100100100001000;
		8'd109: 64'b0100100010000100000010010010000001000000111000010000001100000111;
		8'd110: 64'b0010001000001010010000001010000001100100000111010101000001100000;
		8'd111: 64'b0011000010110100100010010000000001101010000010101000101000100000;
		8'd112: 64'b1101000001010000011100000001000000010000000001001110001000010000;
		8'd113: 64'b1001010000001000011000001000000010000010000001000001000100000000;
		8'd114: 64'b0101001000000010001100000010000000001100010101001101001001010010;
		8'd115: 64'b0010100000000101001001010010111100100001000000000010001010001111;
		8'd116: 64'b0000100000001001001101000001000111011000000000001001000100001001;
		8'd117: 64'b0000101100100011001000000010010100000100011001000000000001110011;
		8'd118: 64'b1010010100000000000001000110011000000100010000000010000000000100;
		8'd119: 64'b0000011001100100011000010000001110000011001011001100000000000010;
		8'd120: 64'b0011001010011001010101000000000011000000000100010000010000101010;
		8'd121: 64'b0000101001110100001110000000000101011000010100000000100100110000;
		8'd122: 64'b0000000100000000000110000000000010000001101110011001000000000010;
		8'd123: 64'b0000001000000000001000100000000000101010000000100000000000000000;
		8'd124: 64'b1100000001000100101001000001000011000100010001100000001010001011;
		8'd125: 64'b0001000010010010000000000000010010000000010000000000000000100000;
		8'd126: 64'b0000010000000011000100010001000000110110010001101000010000001000;
		8'd127: 64'b0100001000000110100000000010000000000010001100010000000000100010;
		8'd128: 64'b0100000000111000000111111001000001100110100010101100000101100101;
		8'd129: 64'b0001001110000010001000001100010100100000001001010010001101000000;
		8'd130: 64'b0000000101000101011010010000100000100001100001000101000100100000;
		8'd131: 64'b1000000000100000001001001000100010000000000001100100000100010000;
		8'd132: 64'b1110000010010010000010000110000010000000000000010000010000000110;
		8'd133: 64'b0100001010000001000100000001110000001001100001010001000000000110;
		8'd134: 64'b0011000000101001010001010001000000010010001001110000101001001100;
		8'd135: 64'b1100000000000000000000000100000000010000001001001011010011010000;
		8'd136: 64'b0000001100010000100010010000110010001010000001000000000010010101;
		8'd137: 64'b0000100100100010000000001001000001011000100110000000100100011000;
		8'd138: 64'b0011001100000100000000000100100000100001000011100000000100000100;
		8'd139: 64'b1000100000000100000001001000010010000101001000000010000101000100;
		8'd140: 64'b0011000010100100100100000100000000000000000000001100000000100000;
		8'd141: 64'b1001010010000001010000100110011011000000010000010000000010000000;
		8'd142: 64'b0000110010001000010010011010100000001000001100000000000000100000;
		8'd143: 64'b0010100000000000100000000011000110000010000000000000000000010100;
		8'd144: 64'b0000000010001001011000000010000010100101001010010001000000000100;
		8'd145: 64'b0100000000000000010011100010000100010001001010100000000000010000;
		8'd146: 64'b0000001000101000010001000000000010000000000000010010010001001000;
		8'd147: 64'b0100000000001000010000100011000011010010100000100000001110100101;
		8'd148: 64'b0000001001000010000000100000000001000001011010000000000000001000;
		8'd149: 64'b0000001101001100000100100100000010100000010010101000010001000001;
		8'd150: 64'b0010101000000110101000010010000010001011000010001010011000100010;
		8'd151: 64'b1010100000000101100001100000110100000000000000111100000000000001;
		8'd152: 64'b1010000000110001000000010000000000000000001000000001000001000000;
		8'd153: 64'b0000001000000000010000100010010010000010100100100001100101001010;
		8'd154: 64'b0000000010100010000101110100000110011011101010100001011000000000;
		8'd155: 64'b0001000110110100000000010010010010110001001101000001001100010000;
		8'd156: 64'b0000000010010010000010000000100000100000100100000000010000000110;
		8'd157: 64'b0010000100000010110010100000000000000000000000000010010010000100;
		8'd158: 64'b0011100000000010010000000000011010100000000101001000001000101010;
		8'd159: 64'b0011000110000110000100001000010010010010101100001000011000001000;
		8'd160: 64'b0000101001000100000010000011101000100000000000000010001000110010;
		8'd161: 64'b0000000000101000110100000010110000000110001001000000000000010000;
		8'd162: 64'b1001001010011000011100000100000001011000101001111000000010000010;
		8'd163: 64'b1000000100000101100000000000100100000001000000000010000100001000;
		8'd164: 64'b1100000100000110000000000000010010000100001011000000000110111100;
		8'd165: 64'b0000000000100110011100010000010100001000101001100000000100010000;
		8'd166: 64'b0000001100010110001100010100000010100001110100010011000001010010;
		8'd167: 64'b1100100000000000100101101001001011000100000000010010011001000010;
		8'd168: 64'b0111000010010001001000100110000000000000000001000000101101000000;
		8'd169: 64'b0010010110101000000000100000001000000001111000011100000000000000;
		8'd170: 64'b0100100000001001000000000011011111000011011110001001110010001010;
		8'd171: 64'b0010000000001011010000000010001100000100101000110001010001101011;
		8'd172: 64'b0001001000001000000000000000100000000000000000000000001000000000;
		8'd173: 64'b0001100000000100011000100000011000000000011000000000101010000100;
		8'd174: 64'b1001000110100010001110100000000100010001101000100001000010010000;
		8'd175: 64'b0101000010010000000000111000100001010000000000000101111010001000;
		8'd176: 64'b0100110001000100000110100001000000000010010110100010010000100101;
		8'd177: 64'b0100000000010101000000100100011010000000000010100011000001001001;
		8'd178: 64'b0100010000100000000101000000001000001000011010100000101100010011;
		8'd179: 64'b0000100101011010000100001010100100000000100010000000000000000010;
		8'd180: 64'b0010001011000000100101010000100000101010000001000100001000010000;
		8'd181: 64'b0010000101000001000000000001100000100000010000000110100010010000;
		8'd182: 64'b0100100100010001000001000000000000000011001110010010000000001101;
		8'd183: 64'b0010001111000000000000010100001000000010101010101000100101011000;
		8'd184: 64'b0000100011101001000010101011100001000000110001000001101000000000;
		8'd185: 64'b0000001101000001010101000001010000000100010100001001001100000000;
		8'd186: 64'b0001000100000010000011001100100000000100001000100010010000100000;
		8'd187: 64'b0000011110000000111100011000000000000001010000000000000000101010;
		8'd188: 64'b1001010010001010101000000001101000001000000000101010100100000101;
		8'd189: 64'b1010000000100000000000000000000000110000011001000000101011000100;
		8'd190: 64'b0000000100000001000000000001001000001001000011010000100010010000;
		8'd191: 64'b0001100001001000001001000111000000100011110011000000100101100110;
		8'd192: 64'b0100000000000001000001010110000011000110010000010001000001000000;
		8'd193: 64'b1100000001001011101010001000000011011101100000010000001000010110;
		8'd194: 64'b0100000010000100000101111000000001000011110001000010001000100001;
		8'd195: 64'b0100001110100000010000000100001011000011001000010100010000010000;
		8'd196: 64'b0100111000000000000101000001010100001000000001000010000100010110;
		8'd197: 64'b0010000001001101000000111001000001010000010000101001100100001010;
		8'd198: 64'b0000000001000000100001100001000101100000000010010001000000000000;
		8'd199: 64'b0000001011011011000010000110000010100100100100011100000010001100;
		8'd200: 64'b0001011000100100000001000000110110001000100101000000011100001000;
		8'd201: 64'b1000001110110000001000110000110000110000001001000011001000001011;
		8'd202: 64'b0000000000000100100000011000010100000000000000100000000010000000;
		8'd203: 64'b0000000010101100010100010000100000001000000111110001001001000000;
		8'd204: 64'b0000000110000000100001000010010010100001000000101010000000100010;
		8'd205: 64'b1001001010010000000000000000010011110000000100000000000100010100;
		8'd206: 64'b1000000000000000101011010000100100000000000000000000110001000010;
		8'd207: 64'b0110000000010011100100000111111010000000001100000101001101000011;
		8'd208: 64'b0100000000001000010000100000000001100000000000000100000001000000;
		8'd209: 64'b0110100000000100101000010010100000000000000010101010100110001000;
		8'd210: 64'b0001001100000001000110000010110101100010001001001000010000100000;
		8'd211: 64'b1011000000000000000001010110100000110000000000000010100001001100;
		8'd212: 64'b0000011110000000000000010110100001010100000000000100000001000000;
		8'd213: 64'b1001000000110000001000000110000010100011000000011001100001010100;
		8'd214: 64'b0001001111000000100000100001000000000110000000001000001100011000;
		8'd215: 64'b1010001001000000000010100000000100000000100000111000000110110000;
		8'd216: 64'b0001001000000000100001000000000000000010000000010001101000000100;
		8'd217: 64'b0111000001000000000100000010000000010000000000000011000001000001;
		8'd218: 64'b0010001000011000010000011010000000000000100100000000100111010001;
		8'd219: 64'b0010000000011000000000010000000000100001011100010100000000001000;
		8'd220: 64'b0001001000000010001100001000011100110001010000000000000110001100;
		8'd221: 64'b0000001010010000100100000000000010010011101000001000000101001001;
		8'd222: 64'b1000001000000000111110010010000100110100000100000000010000111111;
		8'd223: 64'b0000100010000100000000011100000000001001000100010100000011000000;
		8'd224: 64'b1000001000011100000010100010001011011000110000011000110001001010;
		8'd225: 64'b0000001000001000101000000000010010000100000000000101100000100100;
		8'd226: 64'b0110000001000000000010100100000001100001010000000001000011000100;
		8'd227: 64'b0000000011100000000100000010000000100101000000000000100000001001;
		8'd228: 64'b0000000000001000110000010101100011000100110001101000000000011100;
		8'd229: 64'b0000100000010000000010000001000000000000110100000001100100000000;
		8'd230: 64'b0000010100000100000000010000100000000101100000001110111001000000;
		8'd231: 64'b0000111100000000100001010000001010000010000100010000000010000000;
		8'd232: 64'b0000001010000010100001010000000000000000010100100000000001000100;
		8'd233: 64'b0110010100000010000000001000000000011101000010100101000001011100;
		8'd234: 64'b1001001000010011000000000010000000110100000000110100100100110001;
		8'd235: 64'b0100100100001000010100100000001001010000000100010000001010000000;
		8'd236: 64'b0000001001000000000100000010100000100100000001010000101100010000;
		8'd237: 64'b1010101011000000000000000000001100001000010001100100010000000000;
		8'd238: 64'b0100010000100000001000000001000000100111001010000110000000011000;
		8'd239: 64'b0100010010110010001100000000000100000001000100000000000000001101;
		8'd240: 64'b0000001000000000010100010101100100000000101000000000000001101001;
		8'd241: 64'b1000000001000100001001000001011000001000110001000000010000000100;
		8'd242: 64'b0010101010110000110001111000011100100010100010000000000000000001;
		8'd243: 64'b1011010000000101000010000001100011101000111000100000000000000000;
		8'd244: 64'b0100000100000110000000000100010100100010100000100000100010000000;
		8'd245: 64'b0010000000000100000010000001001010110100010000011011100010001000;
		8'd246: 64'b0100000100000100010000000000010000101000000000010000110010100000;
		8'd247: 64'b1100000000010001010100010000000100000001000000000000100000000001;
		8'd248: 64'b0000000001100101011110100000101000010000001010010000000000000001;
		8'd249: 64'b1110000111000110000000000010000010001000000000100100000000011000;
		8'd250: 64'b0100100100100000111001000000010010001000000000001000000000000000;
		8'd251: 64'b0101000010001100000000000101011000000000100100000010000000010100;
		8'd252: 64'b0011001000000010111000000000000000011000000100000011000000000101;
		8'd253: 64'b1000001000010001100000000100100000000000000001000000100010110000;
		8'd254: 64'b0100100001110000010000100010000010010000101000000001000001101000;
		8'd255: 64'b0000000010000001000100010001100001000000000000010100000101100100;
	endcase;
	return out;
endfunction
function Bit#(256) get_msg_bit_page3(UInt#(5) counter);
	Bit#(256) out = case(counter)
		5'd0: 256'b0101101000100000010110001000001001111010110110100100100100011001001010110110001001001111111010111000100101000000001100000110010101111100110011000000011111000101000111001100100001111111001010010111001111000111000001010111100010110101001011001011010101001100;
		5'd1: 256'b0001000101011010100110111011010101011100001001100000100001110010110010011110101111000001110000010100000110100110000101111111100001111101101100101010100010101110111110111111100000000110111010000101100010000001100000110101011010011000010110001101000111000110;
		5'd2: 256'b1001000111100010101000100100000111111111100001111101110011101011001101010111000000011111101111110100101111001111100110100000100101111101000011110010111100000101110011111000100111000010000001011111000001010101001010010001001000111110000000001101101110110010;
		5'd3: 256'b1100101001111110111111011110001010111101000100011000010111010011101001111111111010000100111101011111101111101000101010100001001110001001110100100001001011010110111001001011111011011001001000100111011001101011111001111100011100001100110101111011001001100100;
		5'd4: 256'b0110000010110001111010010111101001000101110000000101001011110111010010010101011001111110100010100110010101000000111001100110010001010010101011111011011110011000100110010000010110101011111000010000001000000101011011101111110010000110101000100011010001001000;
		5'd5: 256'b1111111110011010011000101100110010111011111011110100001011100111001111101110011000000101001011001110100111111011000000101001101101000011110011001000010110111001100010011011110101011100111111001111000100100111001110100001000001011111010001011011101101110010;
		5'd6: 256'b0100101011011101110111011011100101101000111000000111100010011111011111011110000101101101011001110011110110011001111010010000001010110011110001100110011001101011011110010000101000011110101101011111111001111000000110111011110011010110001111110010111111001010;
		5'd7: 256'b1011101011111000110101011111010110100111110000111000100100100000000111100111111101111111111011011011001001000100101010011100101101100010111101111101000111111100010011110111111001001101111111011101000010000010101111011101111011100111100010100010100010110110;
		5'd8: 256'b0111001011101101110010010010011001010100001000000010000110101000100011000101101010101111000110101001101000001111000100000011100010111000110001110000001000010100100110000000100110010010100111000011110001011001000110001010011001000011101010011100110011110111;
		5'd9: 256'b0001011000101110100010000001101010110101000100110100111000100101010001000000011111111010101110110011000011010010111101001111110101101011010110101101111011111011111110100010001100011101100110101001111100111001000000101111110110011000101110100000000011110100;
		5'd10: 256'b1011000101111000110000000010101010111110100000111111111011111000110010100111111110111110001010110100111100101101110011011001101010110011010011000010110110101110001100100111011001101010011100111011010010001111011000000110010100000111101001110101011111111000;
		5'd11: 256'b1001110000101101001011011001100000011010110101001110110110110010110110111101110001100010110000110110000110000001111111101101011110001011110011011101000101000001110100100000010110111000010111010010000010100111101110010111100110100000110000010101000101101100;
		5'd12: 256'b1011101001100000000000100000010111001111110110101001110010101100111001101110111101101001011010010111110001100110101100011111001110101100110001010101001111010001110000110111100100100011001101111100001111101101110110001100000101111100100000000101000010100001;
		5'd13: 256'b1001100000100010001100101011100110000100010011100001111000101110010010111001001000101001010001111110011110100011111110100000001001100100110111111100011100100111110000101100011001101110011101110001110110110010000011100011111100100001111000100000111010110000;
		5'd14: 256'b0001101001110011101001110010100001111010110000000000101000100001011010000110011110001011010011101011011101100111111000000010000011010110100111100110001010100010111111101001110000111001001101110100111101111010101011110010011101010010011110000101101101000110;
		5'd15: 256'b0011011010111111001100010110101110010111111111001000000001001101111111101101011001110110011101100011011110001011110010101011001111001100100100011100010101111111011110101110110111000110100011101111011011011011011000110011010101000110001001010011000100100100;
		5'd16: 256'b0000100110100101110010011101101011000111011000011000010101110101010001111100100011110100101110011111001011111101100010110001000110111011110111100101110100101110111100011111111010000000011111111001001110000011111111100000001010001110100011101100010001110011;
		5'd17: 256'b1011110000011001100101111010101110001000110110001001111001001100111010110011001000110101111100000010111001001100010101011111001000011110000111000011111000000001101011011101000000111010000000111001100000101101110111110010111101000001100001111110101111110101;
		5'd18: 256'b1010001011100100011000110111011111110111100010100001001001001111001010101111001101110101000011001001101001100101111011010001010110110010101011101110010000000101111001001000011110111101111000110000000010000110101111110000010100010001100010001000100000110111;
		5'd19: 256'b0010101110110000000011011101101101001010000101100100001101110101010101011001011011010000011111001001111000111101110110011011100001011111011101110010101110101100011001111010101111101101011111110000110111110100100100110100011000001011000011101111010110001101;
		5'd20: 256'b1010110101001101000111101100000111100100011110100100010101110100011101001101111110110101000000010101111110001001101110010111100011010011010000101110000001100101110010101011000111110110011001010001011111110110000000001000011100010000101111110001011010111001;
		5'd21: 256'b0100101011011010011111100100011101001000010101011011000010001011001100101110110100100011111101011100011100111001000100111110111101000011011001100000010100000111101111100110100110000010001101110111101010100001111000011100010101111011010100001101101100010101;
		5'd22: 256'b0101000011110001110010100000001100010100110110000111010110100000001011111010101000100011100000001101001111011100000100010101111110011100110001111101111100110010100000011101000111111001001111100011101000110001000111110100110101110110111011100000001000111010;
		5'd23: 256'b1111010011011010010110101101011010110011000111011110100100110011100010000110011101011000011001011101101100000101110101101101101011110100111011110111010010000100010001110100100100111100010100110011001100000101111001111111001001111100101011000001011000100110;
	endcase;
	return out;
endfunction
function Bit#(64) get_prev_enc_page3(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1101111011001011010000101100000000011110100100100001110001000000;
		8'd1: 64'b0010111010011100101010001000000011111000011100100000100011000000;
		8'd2: 64'b0000000000000010011001000111010001000000011110110010101000011101;
		8'd3: 64'b0011011011110011000101101001001000111001110111100010001110111001;
		8'd4: 64'b0101000000010001000111110010000011010000001000010000001111101000;
		8'd5: 64'b0000101010111000000010001100011000010000101100101000010011100001;
		8'd6: 64'b0001110011010101001001011100000110111100100001000001000101010001;
		8'd7: 64'b0010011111010100010011100001000000010001100110010101100111010000;
		8'd8: 64'b0101010000100011000000110110100101111100011100010001101000000010;
		8'd9: 64'b0100011000000110101000001000000101000000000001111000100010000100;
		8'd10: 64'b0111000100011000101101001101011010010100000011010011100000001100;
		8'd11: 64'b1001011001110001000010000011000000110001010100111111100100011111;
		8'd12: 64'b1010010001010101110000000100100000000111101100000111010001111010;
		8'd13: 64'b0000110011000010101000000001101000101111110010010011100110011010;
		8'd14: 64'b0101101000010110100010000100000011111100001000110010001000100101;
		8'd15: 64'b0110110000000001000101000000001111010110100001100110010011001001;
		8'd16: 64'b0010010011101110000000010011001011100100101111001101101000010001;
		8'd17: 64'b1110101100000010101001000101001100101000100001100011000001000000;
		8'd18: 64'b1010000110000000101111100000000000110010000010001000011000101000;
		8'd19: 64'b0101101010110111000111111100000010011010110100111001110010000000;
		8'd20: 64'b1010001000001001101000100101101100001001010001111001111111011010;
		8'd21: 64'b0011110111111000100011101011001111101111011100111010101010101101;
		8'd22: 64'b0000000001111010001001100110110001101000001010000000000001000001;
		8'd23: 64'b0011110010011000100000111010110010111101100010010010000110111000;
		8'd24: 64'b1000010110111110110100011011101000000101101001001000100110010111;
		8'd25: 64'b1010101010010101111010111111011110001111001100101110000101100101;
		8'd26: 64'b0001001010011101000001010000100101001011110001011000010010001111;
		8'd27: 64'b0010010110000101000000010000000000100001100000100100101101000010;
		8'd28: 64'b0100101100000010000100100000011110000011011110100000001110000110;
		8'd29: 64'b0110000011100001010100000010100010100001010011010111000110110000;
		8'd30: 64'b0100010010000001001100100000101110010000000001010000110001101000;
		8'd31: 64'b0001000100100010111000011110000101011000101001101100001011000000;
		8'd32: 64'b0100000101010000111000001001100010010000001110000000000000001000;
		8'd33: 64'b1001000001010101011001000110011000000100010101011110101100100000;
		8'd34: 64'b1001010100101010010000010110110100011010100101101100000001101111;
		8'd35: 64'b1010101111011010100001001000100110010000101011101000011110010001;
		8'd36: 64'b1101001101000010101101011111011110001011010010000100111001110101;
		8'd37: 64'b1110011110000001000111110001110001101011110000100001000010000101;
		8'd38: 64'b1000101001000101101101001101011001000100010011000010000000010110;
		8'd39: 64'b0011101110001100110011110001000100110011100010001101100000000001;
		8'd40: 64'b0110010100000110000011100111110011100000110001010100010011001100;
		8'd41: 64'b0011010101010100100110110011000000000100010010001001110000000010;
		8'd42: 64'b1000110101011010010001100001100000000010000100110110010100100010;
		8'd43: 64'b1001101110000101010010011111010010111000000001000101000101001100;
		8'd44: 64'b0101011000011101101101100001110001000111110100010001011101010110;
		8'd45: 64'b0010101110100001110011001001111100000011101100011100000010110011;
		8'd46: 64'b0000110100000100001000100000000100000100001000010100001111000000;
		8'd47: 64'b1110101100011101011011100100000000000000101001000110101011110100;
		8'd48: 64'b0011000000100001011100110001110011111000110010011110001111011001;
		8'd49: 64'b1100001110000011111010100001000001000010100100110000011100010101;
		8'd50: 64'b0000000110001111001000010100111100001101100101010011000100110010;
		8'd51: 64'b1010111010000011001011011000010010111101111000111010010001001110;
		8'd52: 64'b0111010001011010000101010010000110010110000001011100111110010000;
		8'd53: 64'b0101000100010100011101010000000000010000000010000011101001110000;
		8'd54: 64'b0100000111110111010000110101000001111011110111011010010001110001;
		8'd55: 64'b0010011011000111111000001111001000000100100000101100010010010000;
		8'd56: 64'b0100011100000001011111000001000001010000000111000101010011000001;
		8'd57: 64'b0110001000101100011001010110001101000010000111011100110001011100;
		8'd58: 64'b1000000001100011001000110000010001000011010101010110101001001101;
		8'd59: 64'b1000000000111000000110100101001001001100001010010011011101010011;
		8'd60: 64'b1001110110100101001001101010010111000111000000000010000110110101;
		8'd61: 64'b1000100100100001010101000111001011011111111001110101111100100101;
		8'd62: 64'b0110111011000110101001101000000001110010000001001111001101010000;
		8'd63: 64'b1000110010110100001001111011100001001100011000000011010011000000;
		8'd64: 64'b0100010101000011110010000001000100001101111100011100110000010011;
		8'd65: 64'b0110000101011000000110001111100110110000010101001000000010111001;
		8'd66: 64'b0101010000011010000000110001000000011000000010100011010101001110;
		8'd67: 64'b0000011100010101000111100101000001000110010101011010100010010110;
		8'd68: 64'b1000100001100010010001101111110011100111000101100100001001011000;
		8'd69: 64'b1000010000100110000100100010001000100110001101100010100100010010;
		8'd70: 64'b0000000001000000101101000010000110010100010101010100110000101000;
		8'd71: 64'b1011000110111100010110110001011010010111010011100101101100010100;
		8'd72: 64'b1010000100110111011000001001011010000000000100001100001010001010;
		8'd73: 64'b0000110011000100010011000100111100010100000000000001010011000000;
		8'd74: 64'b0111100001101000010000101000000100011110011000011101100101000011;
		8'd75: 64'b0001110010011100000001111110100001000000100111001000000010011000;
		8'd76: 64'b1000010001000010100101110001010100001101000111110001111000000001;
		8'd77: 64'b0100000100000010100010001100001100010100001111010010001111101000;
		8'd78: 64'b1010011011101110000001010101111100010000010010101110110000001011;
		8'd79: 64'b0101100000001111010010111010101001100000100011000000011000111011;
		8'd80: 64'b1110010100010101000001110111010001011000000100011100011101001101;
		8'd81: 64'b1101101010100100001000001000101010111100000001110010010110000001;
		8'd82: 64'b1100100100000000001100000000101000001100101000110111101100100010;
		8'd83: 64'b0010101100100101100101010110010101110011110001010001101101000000;
		8'd84: 64'b0011001010001000100000101110010110000010100001110011111001101000;
		8'd85: 64'b0001011100010001000001100101100000000101110001100011011100000000;
		8'd86: 64'b0011001101100000010011110000011010000010110101100000010101010101;
		8'd87: 64'b0001000011010011100100011001000000010001000110010001010000110101;
		8'd88: 64'b1000111011011010000010010100011110000110001010110000010101000000;
		8'd89: 64'b0011000000100101011000111010011110100011000000010100000100001010;
		8'd90: 64'b1101000001000110000010101000110111110000100111110011001100001111;
		8'd91: 64'b0001100000100110000110000010010100011001000000000001000010010011;
		8'd92: 64'b0000100110111010000010001101101000001011110010100010101010011010;
		8'd93: 64'b0100000110010011011010010001100101101000010100010000101011111010;
		8'd94: 64'b0010101000000101001010000111100001100010100001000000101101001000;
		8'd95: 64'b1100000101110001101100001000010001100000010001011111010000100100;
		8'd96: 64'b0010001110101001010110110010101100000000100001010010010111101100;
		8'd97: 64'b1001111100101000001110101011000010100001001010101111100000000101;
		8'd98: 64'b0010000000000010101000110001001101110011001100100100010000100010;
		8'd99: 64'b0111100111000110001000001101000110010000001001001110010011000000;
		8'd100: 64'b1001111100001001111100011000100111011101001000001101000110100100;
		8'd101: 64'b0011100100100000010000001110011101011000000001100100010100010100;
		8'd102: 64'b0101000011010110011110100101011101111000101001001100100000000110;
		8'd103: 64'b0101010101000011001010001010000010000011001000100110001000010010;
		8'd104: 64'b0000111100000001000100000000111110010010010010111111110001011011;
		8'd105: 64'b0010001000000111011101010000111000000000000000110010010000010010;
		8'd106: 64'b0000111100110000001010001001000000100111001100110000000011010001;
		8'd107: 64'b1001110010100001010001110001100010010001000010000000001001100000;
		8'd108: 64'b1001011100001000001100110010011000011001000011011110101100111000;
		8'd109: 64'b0100101010100100000010110010000011001010111000110100011100100111;
		8'd110: 64'b0110001000101011010000001010010001100100000111010101010001100100;
		8'd111: 64'b0011000010110100100010010001001011111010101011101000101101110000;
		8'd112: 64'b1101000001010011011100000011010000010000100101001110101000010000;
		8'd113: 64'b1001011000001000011111001000000010000010000011000011000110000000;
		8'd114: 64'b0101001000001010001100000010000000001101010101011111011001010011;
		8'd115: 64'b0010100000100101001101111110111100100001010001000010011111001111;
		8'd116: 64'b0000100110101001001101000001100111011001000001011011011100001001;
		8'd117: 64'b0111101100100011001010100010010101000100011001110000000001110011;
		8'd118: 64'b1010110100000010001011000111011001000110110010100010010000000100;
		8'd119: 64'b0000011101100100011000111000001110010111001011001101010000000010;
		8'd120: 64'b0011001011011111010101000000000111000010000110010000010001111010;
		8'd121: 64'b0100101111110111001110100000001111011100010110000000100100110001;
		8'd122: 64'b0000010110010101000110100000001010000011101110011001100101001011;
		8'd123: 64'b0011001001000000001100100000000000101010010000100000101100000000;
		8'd124: 64'b1100101001000100101001100001010011000100011001100010101011101011;
		8'd125: 64'b1011000010010010101000000100010010000000110000101001010010110000;
		8'd126: 64'b0110010001001011000101110001000000110110010001101001010000001010;
		8'd127: 64'b0110001010110110100000000010010100100010001101010100000000100110;
		8'd128: 64'b1100110000111010000111111111010001100110100010101100010111101101;
		8'd129: 64'b0001101111000111101000001110011111100000001001011110001101000010;
		8'd130: 64'b0100000111000111011011010000110100111001100001010101000111100111;
		8'd131: 64'b1000000000100010011001101000100010000000001011101100000100010000;
		8'd132: 64'b1110000010111011010010100110000010000100000000111000110001000110;
		8'd133: 64'b0100001010000001100110000001110100001011100101010101011111000110;
		8'd134: 64'b0011001000111011010001010101110100010010011001110000111001001100;
		8'd135: 64'b1100101000100100010100000100000100011000101001001111110111010000;
		8'd136: 64'b0001011100110000101110110000111011001011000111001010010110111111;
		8'd137: 64'b0000100100100111000000111001100001011001101110000000100100111000;
		8'd138: 64'b0011001100000100000000001100100000111001001011100010000100011100;
		8'd139: 64'b1001110000000110100011001000010110001101001001010010110101010100;
		8'd140: 64'b0011001010101100100100000100000100001000000000101100101011100011;
		8'd141: 64'b1001010010000001010000100110011011010110110000010000101010000100;
		8'd142: 64'b0100110010101000111110011010100000001000001111000000000000101000;
		8'd143: 64'b0010101000011000100000000011001110110011000000100000000000010111;
		8'd144: 64'b0000000010001001011001100110000010100101011110010001001000010100;
		8'd145: 64'b0100001000011000011011100011000100110001001010100110100001010000;
		8'd146: 64'b0000001000111101010001001000000111000000100010110011010001001111;
		8'd147: 64'b0110001001001000010010100011001111010010100011110100001110110101;
		8'd148: 64'b1100001101000010010000100000000001000001011010000000010000001001;
		8'd149: 64'b0010101101001110000100100110011110100111011011101000010001001111;
		8'd150: 64'b0010101010011110101100110110010010011011100010001010011000100010;
		8'd151: 64'b1010100000000101101001100000110110101010000010111100000100000001;
		8'd152: 64'b1110000000111011010001010011101000010101001101001001000001101010;
		8'd153: 64'b0000001000001000010100110010010010000011110110100001100101001010;
		8'd154: 64'b0001101110101010000101111111010110011111101111110001011010001000;
		8'd155: 64'b0001101110110110000001110011010011111011101101000001011100010101;
		8'd156: 64'b0000010010010010000110110000100000101000110100000000110000000110;
		8'd157: 64'b0010001100000010110010101000000010000000000000000010010010000100;
		8'd158: 64'b0011100000010010010001000100111010100010001101101000011000101011;
		8'd159: 64'b1111010110010110110100101000011110010110101101101000011000101000;
		8'd160: 64'b0011101101011110010010010111101001100000101000100110001011111011;
		8'd161: 64'b0001000000101000110100000010110010000110001011100001000000011000;
		8'd162: 64'b1011001110011001011101000100000001111000111001111110001010000011;
		8'd163: 64'b1000000100000101100110010000100101000001000000010010000100001000;
		8'd164: 64'b1101000100000110000100100000010010100100001011000000100110111100;
		8'd165: 64'b0000000000110110011101010010010100011000101011101001000100010010;
		8'd166: 64'b0000001100010110001100110111000010100101110111010011100101010111;
		8'd167: 64'b1101100001000000100101101001001111000100100000010110011001000010;
		8'd168: 64'b0111001010010001001000111110000000000001111001000100101101010011;
		8'd169: 64'b0010010110101010000110110000001000000001111001111100110000011010;
		8'd170: 64'b0110110000101101000000001011111111100111011110001001111010001010;
		8'd171: 64'b0010000000001011111000000010001101110100101000111001010011101011;
		8'd172: 64'b0001001000001010000000000110100100000100000000000001001000001000;
		8'd173: 64'b0001100100000100011010101011011000000010011000000000101010100110;
		8'd174: 64'b1001000110110110001110100000000100011001101001100101110011010001;
		8'd175: 64'b0101000010010000010000111000100001010000100000000101111010001000;
		8'd176: 64'b0100111101010100000110100011000100000010010110100110010000110101;
		8'd177: 64'b0100000001010101000001100100011110001000000010110011010001001001;
		8'd178: 64'b0100011000100000000111010110001001001000011010110000101101011011;
		8'd179: 64'b1000100101011010010110001010100100000000100110100000001000000110;
		8'd180: 64'b0010001011000000100101010000100000101010000101011111001101010100;
		8'd181: 64'b0010000101000001100000000001110000111000010001110110100010010000;
		8'd182: 64'b0100111101011001100001000001100100010011001110010010010000111101;
		8'd183: 64'b0010001111001000000000010100001001100010101010101110111101011000;
		8'd184: 64'b0100100011111001000110101011101001000001111001100011101110000000;
		8'd185: 64'b0001001101011001110101100001110000000110011101011001001100010001;
		8'd186: 64'b0001010101000010001011101100100000000100011000100010010100100100;
		8'd187: 64'b0001011110010000111110011001000100001001010110000000000100111010;
		8'd188: 64'b1011011010001010101010001001101000101010101001101011100110010111;
		8'd189: 64'b1110000101100000001000110100010001110001011001000100101111100100;
		8'd190: 64'b0100000100000001000100000001011100001001000011010100101010010010;
		8'd191: 64'b0001100101001000001001000111100101100011110011000100100101100110;
		8'd192: 64'b0100000001100001000011010110000111010110010000010001000001100000;
		8'd193: 64'b1100011001001011111010011001010011111111100000010000001101010111;
		8'd194: 64'b1110000010000100010101111001000001010011110001001011001000100001;
		8'd195: 64'b0101001110100010010001100111001011000011001100011101010000010010;
		8'd196: 64'b1110111010100100010101101011011100001110000001010010010101010110;
		8'd197: 64'b0111000001001101001010111001100101111000010110111001101100001110;
		8'd198: 64'b0000000001001101100011100001000101100010000010010011100000000000;
		8'd199: 64'b1010001011011011000010001110000010110100100100011100100010011100;
		8'd200: 64'b0001011000100100110101000010110111001000101111000100011100101001;
		8'd201: 64'b1000101110110010001000110010110100110010001101000011001000101011;
		8'd202: 64'b0000001000100100100000011100010111000000100000101010000110000000;
		8'd203: 64'b1000000110101101110110010010110000001000000111110001101001001010;
		8'd204: 64'b1000000110010110100001000010010010100011000000101010001000100010;
		8'd205: 64'b1001011011010000010001110000010011110110110100000100000100011101;
		8'd206: 64'b1100100000101000101011010100100100000010101001000000110001100110;
		8'd207: 64'b0110010101010011100100000111111010010000101100110111001101010011;
		8'd208: 64'b0101000000101000010000100011000001100000000010100100000001000100;
		8'd209: 64'b0110100000000111101000010010100001100000000010101010100110011000;
		8'd210: 64'b0001001100000011010110010010110101110010011001001001010100100000;
		8'd211: 64'b1011000000110000001001010110110100110000010010000010110101001100;
		8'd212: 64'b0000011111000000000110010110100001010101001000010100000001000110;
		8'd213: 64'b1011000000110001011000000110010010110011000000011001101001010100;
		8'd214: 64'b1001111111000000100100110001110100010110010000001010101100111100;
		8'd215: 64'b1110001111000000000010110000001110000001100000111000000110110001;
		8'd216: 64'b0111001000000101110001100000000100000010000010111001101001000110;
		8'd217: 64'b0111000001000000000100000010000000010011010000000011010001000001;
		8'd218: 64'b0010001011011000011000011010011010000001110100000010100111010001;
		8'd219: 64'b0010000000011000100100010011000100100101011100010100011100011000;
		8'd220: 64'b0101001000001110101101011000011101110011010101000010000110001100;
		8'd221: 64'b0000001111111000101100110001000010010011101110001000000101001001;
		8'd222: 64'b1000011000100000111111010010010100111100100100000000110000111111;
		8'd223: 64'b0000101110000111001001111100000011001001100100010100000011100000;
		8'd224: 64'b1000011010011100000010101110001011011100110000011000110001101010;
		8'd225: 64'b1010101000101001101000000000110010100100001010011101100000101100;
		8'd226: 64'b0110000101000100010110101100000101100001010000000001000111100100;
		8'd227: 64'b0010011011100000000101010010110101111101001000000010101100001001;
		8'd228: 64'b0000000000001000110000110101100011000100110011101000101100011100;
		8'd229: 64'b0100100000011000010010010101001000110001110101000001100100000100;
		8'd230: 64'b0100111111000100101000110001100000000101110000011110111001010001;
		8'd231: 64'b1000111100010000110001010100001010000011010100011000010010000000;
		8'd232: 64'b0000001010000010100101010010010000000010010100100000010001010101;
		8'd233: 64'b1110011101000010000000001000001001011111001010100111000001011100;
		8'd234: 64'b1011011010010011000010001010000000110100100100111110100100110011;
		8'd235: 64'b0110100100111000010110100001001101110100000100010011001010000100;
		8'd236: 64'b0000001001000001100100101010100000100100000001010100101100011000;
		8'd237: 64'b1010111011010111001011011000001100001011110001101101011000010100;
		8'd238: 64'b1100011011100000001000000001100101100111001111000110110000011000;
		8'd239: 64'b0101011010110011101100000000100110100001001100000000000000111111;
		8'd240: 64'b0110101000000010010100010101100100000010111010000000000111101001;
		8'd241: 64'b1110001001000100101001000001011010001000110011011010010000011100;
		8'd242: 64'b0010101010110000110001111100011110100010110010001000010011001001;
		8'd243: 64'b1011010000010101000010000001100011101000111001110001010010010000;
		8'd244: 64'b0100101101000110000000001100010100100011100001100000101010011010;
		8'd245: 64'b0010000010100100000010010011001010110100110000011011100010001000;
		8'd246: 64'b0100110100001100010000000000010000101100001000110000110010111010;
		8'd247: 64'b1100100100010001010110110010000100000001010010000010100000110001;
		8'd248: 64'b1100000001100101011110100000101001010001101010010010100001001001;
		8'd249: 64'b1110000111010110000001000010000011001000000000100100011000011011;
		8'd250: 64'b0111100100101110111001100001111110001001000010001001010000000100;
		8'd251: 64'b0101000010001100000101100101011000001100110111110111110000010110;
		8'd252: 64'b1011001000000010111000001000010101011010000100000011100010000101;
		8'd253: 64'b1000001000010001100010010100110000010001001001000001100011110100;
		8'd254: 64'b0111101111110000011010100011000010010000111110010001000101111000;
		8'd255: 64'b0000000010000001000100010001100001000001000100010101010101100101;
	endcase;
	return out;
endfunction
function Bit#(256) get_msg_bit_page4(UInt#(4) counter);
	Bit#(256) out = case(counter)
		4'd0: 256'b1001111010001100001111010101001101010100010010011100100111101010101010100000111010110001101100100011001010001100001110110001101000011100111011000001100100010101100110100011101101011111000010101110011011101101010100101100111110101111000001101110100000010111;
		4'd1: 256'b1001100100100100000111011100111010110111001000101001011011101100111110011000111011111001111001001011101000000111000001100001111010000111111000011110110000011010111101011010001101110100100001110000010011110010011001110011111000110110101010001100110101110111;
		4'd2: 256'b0101100100101111111001111011100100011100111110111110110001111111010011110000100001101001100111000000101101000100100010010110001000110011000100011011111010110000101100001001111010010111010011001100110010110101111000000010011011001001111100001001000111010110;
		4'd3: 256'b1101101110100100110101111011001101011011111011100101000001100000110010001010101011011001100000000111100100000000111010100001110001000111011110111000111000000101001110001101110111110101000010000100111101100010100110010010100000011001101100101010000110110000;
		4'd4: 256'b1111110101101000000001000100110011011011001100110000100001000011111000001101101100001011001001010111001011001101011010001011110111001100100001001000011101000110000110100010110010101111010011110100110011000000101100101101010110011010101001001101101011111101;
		4'd5: 256'b0000101010000000110010110000011100110101001001110000010101010001101111011011111110101111011110011101001101110001111011011101111100100100111110100110111000010010000111110111100110110111100111001011100001011010010010111000001100000001010110001001000101101010;
		4'd6: 256'b1111010001000011110111101000011011101010101001101011000110101001010111111000110110001110111110011110000011101010110110111000100111010000001100100000111000011011010100111001100000011011011000010101111001111011000101110010000100111011100100110011110011111010;
		4'd7: 256'b1001101111000101110000010011001001011011110111111011110001111001100101010001000111100110000110111100010010111111110101100111111011110101101111101010111011000111001010111000100010100010100011101001001100000010010100010100001000101101101101000011011011010010;
		4'd8: 256'b1110011010100001101100011110101110001000100110111001100100010011101111110011010100000001110100011101001000100101111001100000010110111110110101001000100111110110111110000110110001011000101011011011011111010110001111100000001011100000011110110001000010001100;
		4'd9: 256'b1101000011000110101000011110001111010110111101001110010100010111110101111011001011011000101000111111010010010100010010000110100010011001101011000010011010001100010101101010010101101011111011110010100111100111100011101001101000110111100001100101001111101010;
		4'd10: 256'b0011110111010101110011110100111110001000010101010111011110010011101100101100110000110010001110001111010001011000010101110111001001111000110110110001001010101000111100101000101011000110110100000011000011110001000010011001110110111100111000000101110110101110;
		4'd11: 256'b1111111100000011001110101110110101101001001001100110001011000111001000011101100010000000011001000010001010101001000010011110011011101001111101001011011111110101100011011000010111110101101110001000101101101010000100111011101100001101110000001111101010010100;
		4'd12: 256'b0011010110000100100111000010100111100010110101110110000111011100001111110000001010111101010101111001100110110101011111100110000001101001111010001001110111000111001001000111010010010110011001100101011011111101000011001111101000011110001100000101101101111101;
		4'd13: 256'b0010111101111001010010101000110110100110001100110101100100111010110001011110110000100110110011011101010000110001010001000101011010100001100001110010011101101100100100111001101110110001111110110000101110101101001100001111010101011011011011001011111101100011;
		4'd14: 256'b0100011000011101100000101110011000010110100111110100010110000101110010110110000100001000000100101111011011010010011000100101100011010000010111001001110110010101111001000111100100110101011111100000010011100111011001010010010000111010111011000110011100100011;
		4'd15: 256'b1000101100011111001001010001101011110110001010110101101101000100111110111110001010000011011110100101110010010000110111101100100100111011000111001100111110001101110111100000010111100010000111011100110110110111001010011010010111000100000001001101101100110101;
	endcase;
	return out;
endfunction
function Bit#(64) get_prev_enc_page4(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1111111011011011111101101100000010111110100110111001111011001000;
		8'd1: 64'b0010111010111110101010011010001011111010111100100010100111000010;
		8'd2: 64'b0010010000000010111011100111010001100010011110110110101100011111;
		8'd3: 64'b1011011011110011000101101001001000111001110111100010001110111001;
		8'd4: 64'b1101000001010011000111111110100011010001101000010100101111101000;
		8'd5: 64'b0000101010111000000110011100011000111000101110101000010011100111;
		8'd6: 64'b0101110011010101101001111110000110111100100001010101010101010001;
		8'd7: 64'b1011011111010100011011100001000000110001100110010101101111010001;
		8'd8: 64'b0101011100100011000010110110100101111100111100010101101000000010;
		8'd9: 64'b0101011010000110101110001000001101000010100011111100100010000100;
		8'd10: 64'b1111000110011000101111001101011010110100000011010011100001001100;
		8'd11: 64'b1001111001110001000111000011000000110001011101111111100110011111;
		8'd12: 64'b1010010001010111110001100101100001000111101100001111010101111010;
		8'd13: 64'b0010110011000010101000001001101000101111110010010011100110011010;
		8'd14: 64'b0101101010010110101010000111001011111100011100110110001010100101;
		8'd15: 64'b0110110100000011011101001010001111010111100001101110010011001011;
		8'd16: 64'b0010010011101110000000011111001111100100101111001101101000010001;
		8'd17: 64'b1110101101100011101001000101001110101000100001100011000001000100;
		8'd18: 64'b1010000110001000111111100100000000111010000010001100011000101000;
		8'd19: 64'b0101101010110111101111111100001011011010110100111001110110100001;
		8'd20: 64'b1010101000011101101011101101101101101011010101111011111111011010;
		8'd21: 64'b0011110111111011110011101011001111101111111110111010111110111101;
		8'd22: 64'b0000100001111010001001100110110001101000011110000000000001101001;
		8'd23: 64'b1011110010011000100000111011110110111101101010010010000110111001;
		8'd24: 64'b1000010110111111110100011011111100000101101001101000100111010111;
		8'd25: 64'b1110101010010101111010111111011110001111011101101110000101110101;
		8'd26: 64'b0001001010011101000001011100110101001111110101111000010010011111;
		8'd27: 64'b0010010110011101010000010010000100100101100000100100111111000110;
		8'd28: 64'b0100101100100010100110100000011110100011011110100000001110000110;
		8'd29: 64'b0110011111100001011100000010110010100001010111011111000111110010;
		8'd30: 64'b0100010010000001001100100100101110010000000001010001110001101001;
		8'd31: 64'b0001001100100110111110111110001101111100101001101100011111001100;
		8'd32: 64'b0100000101011000111000001101100010010000011110000001000010011000;
		8'd33: 64'b1001000101010101011001000110011100000100011101011110101100101110;
		8'd34: 64'b1001010110111010110000110110110100011010101101101110000001101111;
		8'd35: 64'b1011101111111011101001101001110110010000101111111001011110010001;
		8'd36: 64'b1101001101010011101101011111111110011011010010110100111001111111;
		8'd37: 64'b1110011111000011010111111101111011101011110000101001001010010101;
		8'd38: 64'b1100101001001101101111001111111001001101010011001010000011010110;
		8'd39: 64'b1011101111001100111111110001000100110011100010001101101100000001;
		8'd40: 64'b0110010100010110000011101111110011100000110111010100010011001100;
		8'd41: 64'b0011010101010100100111110011001000000100010110001001110000000010;
		8'd42: 64'b1000110101011011010001100001101010000010010100110110010100100110;
		8'd43: 64'b1001101110000101110110011111010010111000000101000101000101011100;
		8'd44: 64'b1111011100011101101101111011110001010111110100110011011111010110;
		8'd45: 64'b0010101111110011110011011001111111000011101110011100011111110011;
		8'd46: 64'b0000110100000100001100111101010100000101001000010100001111000100;
		8'd47: 64'b1110101100011101011011100100000011000000101001100110111011110100;
		8'd48: 64'b0011101110100001011111111001110011111000110010111110111111111101;
		8'd49: 64'b1110101110000011111011100011010011000010100100110000011100010111;
		8'd50: 64'b1000100110001111001000110100111100001101101101010011000100110011;
		8'd51: 64'b1010111010100111001011011001011010111101111000111011010001001111;
		8'd52: 64'b0111010001011110100101010010001110010110000001011100111110010011;
		8'd53: 64'b0101000100010100011101010000000000010000100110000011101001110000;
		8'd54: 64'b0101000111110111010100110101100001111011110111011010010001110001;
		8'd55: 64'b0010011011000111111001001111001010000100100001101100010110110010;
		8'd56: 64'b0100011101000101011111000001000111010101100111000101110011011001;
		8'd57: 64'b0110001100111111011101110110011101100010010111111100111001011100;
		8'd58: 64'b1110000001100011001001110000010001000011010101010110111011001101;
		8'd59: 64'b1000010000111000100111110101001011001100101010010011011111010111;
		8'd60: 64'b1001110110100101001001101010010111001111100001000010011110110101;
		8'd61: 64'b1100100100110001110101000111111011011111111101110101111101100101;
		8'd62: 64'b0110111011000110101001101000000001111010000001101111001101010101;
		8'd63: 64'b1000110010110100011101111011110001101100111110000011011011100110;
		8'd64: 64'b0100010111000011110010000001000100001101111111011101110001110011;
		8'd65: 64'b0111100111011000100110001111100110110010010101011000101010111001;
		8'd66: 64'b0101111010011010010000110111001000011000101010100011010111011111;
		8'd67: 64'b1110011100010111000111100101010101100110010101111110110110010110;
		8'd68: 64'b1001100001100010010101101111110011110111000101101100011011011110;
		8'd69: 64'b1100010100111110000100110010001011100111001101100010101100010010;
		8'd70: 64'b0001010111000100101111000111000110011100110101010100110000101000;
		8'd71: 64'b1011111110111101011110110001011011010111010111100101101110111100;
		8'd72: 64'b1010000100110111011000101001011010000001000100001100001010001110;
		8'd73: 64'b0000110111000101111011000100111100011100010000001011010011000100;
		8'd74: 64'b1111100101101001110001111000000110111110111100011111110101011111;
		8'd75: 64'b0001110010011100000111111110100001000000100111001000100010011111;
		8'd76: 64'b1000110001000010100111110011010101111101100111110001111111011001;
		8'd77: 64'b0110010100001010100010001100111100010100001111010010111111101100;
		8'd78: 64'b1010011011101111000001010101111100010001010010101111110100001011;
		8'd79: 64'b0111100000001111110011111011101001100000101011000000011000111011;
		8'd80: 64'b1111010100110101010011110111010101011100010111011100011111101101;
		8'd81: 64'b1101111010100100101000001100101010111100000001111011010110000001;
		8'd82: 64'b1100100101000000001100000000101011001100111000110111101100101010;
		8'd83: 64'b1010101101100111100111010110010101110011110001110001101111000100;
		8'd84: 64'b1011001010001100100001111110011110110110100001111011111011101100;
		8'd85: 64'b0101011100010001100111110111101100000101110001100011011110010000;
		8'd86: 64'b1011001101100000010011110001011111010010111101101100010101110101;
		8'd87: 64'b1001000011010011100110111001000010010001010110010001010110110101;
		8'd88: 64'b1000111011011110000111010101011110000110101011110000110101000001;
		8'd89: 64'b0011101100100101111000111010011110100111001100110100000100011010;
		8'd90: 64'b1111000001000110000010101100110111110100101111110011011100001111;
		8'd91: 64'b0001100000101110000110000011010100011001001000000001000010010111;
		8'd92: 64'b0000100110111010011011001101101000001111110010101010101011011010;
		8'd93: 64'b0100110110011011011010011001100101101001110100110010101111111010;
		8'd94: 64'b0110101110001101001010010111100001111110100001000100111101001000;
		8'd95: 64'b1101010101110001111100101000110011100000110101011111111000100100;
		8'd96: 64'b0010001110101001010110110010101100001001111111010011010111101100;
		8'd97: 64'b1001111110101010111110101011100010100111001010101111110000000101;
		8'd98: 64'b1110001000010011101001110001001101110011001100100110010000100010;
		8'd99: 64'b0111110111100110011000101101000110010001001101001110010011100000;
		8'd100: 64'b1001111100001001111100011000100111011101001100001101000110100100;
		8'd101: 64'b0011100100100000010001001110011101011000001001100100010110010100;
		8'd102: 64'b0101000011011110011110111101011101111100101111001100111001010111;
		8'd103: 64'b0111011101000011001010001010000010010011011000100110001110010010;
		8'd104: 64'b0000111110001001101100010000111111010010010010111111110001111011;
		8'd105: 64'b0010001000000111011101110000111100000101000101110010010100111010;
		8'd106: 64'b0000111110110011001111001001100110101111001100110000011111010001;
		8'd107: 64'b1011110110110001010001110011100010010001000010000010001001100000;
		8'd108: 64'b1111111100101110001100110010011000011111000011011110111100111000;
		8'd109: 64'b0101101010100110000110111011000011001010111001110100011100100111;
		8'd110: 64'b0110011001101111010000001010010101100100001111010111010011100100;
		8'd111: 64'b0111000110110101101010010011001111111011101011101000101101110000;
		8'd112: 64'b1101000001010011011101100011010010010000110101001110101001110100;
		8'd113: 64'b1001011000001110011111001100100010010010000011000011111110000000;
		8'd114: 64'b0101001000001011001100010010000110011101010111011111011001010011;
		8'd115: 64'b0110100000100101001111111110111101100101110001000010111111101111;
		8'd116: 64'b1000110110101011101111010001100111011001000001011011011100101001;
		8'd117: 64'b0111101100101011001010101010010101001100011001110010100011110011;
		8'd118: 64'b1010110111000010001011001111011001000110110011100010010000000100;
		8'd119: 64'b0101011101110100111000111000001111010111011111001101010000000010;
		8'd120: 64'b0011001111011111010101000000000111000010010110110000010001111010;
		8'd121: 64'b0101101111110111001110100000001111011110010111000000100100111001;
		8'd122: 64'b1000010110010101100110100001001010010011111110011001100101001011;
		8'd123: 64'b0011001001010010001100100000000000101010010100100100101101000000;
		8'd124: 64'b1100101001000100101001110001010011001100011011100010101011101011;
		8'd125: 64'b1011000010010011101000001100010010000000110011101001010010110010;
		8'd126: 64'b0111010001001011000101110001101000110110010001101001011000001010;
		8'd127: 64'b0111001010110110100000011010010100100110101101010100000000100111;
		8'd128: 64'b1100110000111010010111111111010001100110110010101100110111101101;
		8'd129: 64'b0111101111000111111011001110011111101010001011111110011101000110;
		8'd130: 64'b1100000111000111011011111000110100111001100001010101110111100111;
		8'd131: 64'b1000000010110010011001101001100011000010101011111100010110010010;
		8'd132: 64'b1110000110111011010010100110001110000101010000111000110001000110;
		8'd133: 64'b0100001010000011100111000101110101001011110101010111111111000111;
		8'd134: 64'b1011001010111011111001010101110100110010011011110001111111011101;
		8'd135: 64'b1100111000110100111100010101000110111000101001001111110111010010;
		8'd136: 64'b0011011100110000101110110001111011001011000111111010110110111111;
		8'd137: 64'b1001100100110111000010111101100101011001101110101100110100111001;
		8'd138: 64'b0011001100100110000000001100110000111001001011100010100100111100;
		8'd139: 64'b1001111000001110100011001000010110001101001011011010110101010100;
		8'd140: 64'b0111101010101100100101000100100100001010010000101100111011100011;
		8'd141: 64'b1001010010000001010100101110011011010110110001010000111010001100;
		8'd142: 64'b1100110010101000111110011010101010011001001111000000000000101010;
		8'd143: 64'b0010101000111010101000000011001110110011010000100010001001010111;
		8'd144: 64'b0000000110001001011001110110100110100111011110010101101100111100;
		8'd145: 64'b0100001000111001011111110011001100110001001010100110100001110010;
		8'd146: 64'b0000101000111111111001001000100111000000100010111011010001001111;
		8'd147: 64'b0111001001001100010010101011101111010010111011110100011110110111;
		8'd148: 64'b1100001101000010010000100000000001011001011010000000010001001101;
		8'd149: 64'b0010111101001111000111100110011110100111111011101000010011001111;
		8'd150: 64'b1010111010011110101101110110011010011011100010001010111000101010;
		8'd151: 64'b1010101000011101101011101000110110101010000011111100000100001001;
		8'd152: 64'b1110000100111011011011011011101000011101001111001101101001101010;
		8'd153: 64'b1000001000001000010100111010011011010011111111100111110101001010;
		8'd154: 64'b0001101110101010100101111111111110011111101111111001111110101000;
		8'd155: 64'b1001101110110111001101111011010011111011101101010001011100010101;
		8'd156: 64'b1000011010010110000110110010110000101010110110000000110100001110;
		8'd157: 64'b0010001110000010110011101000010010010000000001001010110010000100;
		8'd158: 64'b0011110000010011011001100100111110100010001101101010011000101011;
		8'd159: 64'b1111011110110110110100101001011110010110101101101010011000101010;
		8'd160: 64'b0011101101111110010010010111101001110001111000100111001011111011;
		8'd161: 64'b0001100100101000110101000010110010010110001011100001001000011100;
		8'd162: 64'b1011101110111111011101011100001001111100111001111110101010000111;
		8'd163: 64'b1001000100100101100110010000101101000001100000010010100101001001;
		8'd164: 64'b1111100100100111101100110000010010111100001011000000100110111100;
		8'd165: 64'b0000000000110110011101110010010100011000101011101001000100010011;
		8'd166: 64'b0010001101010111001100110111000010100101110111010011110101010111;
		8'd167: 64'b1101100001000000110101101011011111000110110000010110011011000010;
		8'd168: 64'b0111001010110001001000111111000000100101111001000100101101010011;
		8'd169: 64'b1010010110101010000110111010001000000001111001111100110001011010;
		8'd170: 64'b0110110010101111100000001011111111101111111111101001111010001010;
		8'd171: 64'b0010001000101011111000001010101101110101101000111001011111101011;
		8'd172: 64'b0001011000001010000000001110101100100100010110000001001100001000;
		8'd173: 64'b0011100100000100011010111011011000010011011001110010101011100110;
		8'd174: 64'b1101100110111110001110100001000101011001101001100101111011010011;
		8'd175: 64'b0101000010010000010001111000100001011000100000100101111010101010;
		8'd176: 64'b0100111101010110010110100011000101000010010110100110010010110101;
		8'd177: 64'b0100100001010111101001100100011110001100010010111011110001001001;
		8'd178: 64'b0100011001100010000111110110001001001001011010110001101101111011;
		8'd179: 64'b1011100101011010010110001010110100100000110110100100001000000111;
		8'd180: 64'b0010011011000000101101011000100100101010000101011111101101010101;
		8'd181: 64'b0010000101000101110000010101110000111001010001110110100010010000;
		8'd182: 64'b0100111101011001100001000011100100011011011110010010010100111101;
		8'd183: 64'b0011001111101000011000110100101111100011101010101110111101011010;
		8'd184: 64'b0100100111111101000110101011101011001001111001100011101110000010;
		8'd185: 64'b1001001101011001110101101101110100010110011111111011001100010101;
		8'd186: 64'b0001010101000010001111101101100000000100011000101111010101100100;
		8'd187: 64'b0001011110011000111110011001000110011101010110000011000100111011;
		8'd188: 64'b1011111010001010101010001001101010101110101001101011100110010111;
		8'd189: 64'b1110000101100000001110110110010001110001011001000100101111100100;
		8'd190: 64'b0100001101000011000100000001011100001011000011010100101010010010;
		8'd191: 64'b0001100101101100011001000111101101110011110011000110100101110110;
		8'd192: 64'b0100011101100101000011010110000111110110010000110001000111100000;
		8'd193: 64'b1100011001001011111010011011010011111111100010010110001101110111;
		8'd194: 64'b1110101010000100011101111001110101010011110001001011011011110001;
		8'd195: 64'b1101011110100111010001110111011011000011111100011101011010010110;
		8'd196: 64'b1110111010101100010101101011011100111110001001010010010101110110;
		8'd197: 64'b1111000001001101001010111011100111111000010110111001101100011110;
		8'd198: 64'b0000010001001101101011101001000101110010000011010011100000000000;
		8'd199: 64'b1010001011011011000010001110100010111101100111111100100011011100;
		8'd200: 64'b0001011000110100110101000010110111001000101111011100011100101001;
		8'd201: 64'b1010101110111110001100110010110100111010001101000011001000101011;
		8'd202: 64'b0000001110100101110100011101110111001010100001111011000110000100;
		8'd203: 64'b1000101110101111110110010010111100101000100111110001101111001010;
		8'd204: 64'b1000000110110110100001001111110010101011011000101010011000100110;
		8'd205: 64'b1011011011011000011101110001011011110110110101110100000110011101;
		8'd206: 64'b1110100000101010101011011101110100101010111011001000110001101110;
		8'd207: 64'b0110010101010011111110000111111010010001111100110111101101110111;
		8'd208: 64'b0101000000101000010010100011011001101100010110100100000001000110;
		8'd209: 64'b0110100000101111111000010010100001100000100010101010100110111000;
		8'd210: 64'b0001011101000011010111010010110101110111011001101001110101100000;
		8'd211: 64'b1011010000111100001001010111110110110000010110000110111101001100;
		8'd212: 64'b0000011111100000000110011110100011010101011000010100000001000110;
		8'd213: 64'b1011000100110001011111100110010010110011001101011011101001010100;
		8'd214: 64'b1001111111100010100110110101111110010110010011101110101100111110;
		8'd215: 64'b1110001111001100000010110000001111000001100100111000000110110001;
		8'd216: 64'b0111011000000111110001110000010100000110000010111011101001100110;
		8'd217: 64'b1111001001001010011100000010001001010011010000000111010011000001;
		8'd218: 64'b0010001111011001111100011011011010000001110100001110110111010101;
		8'd219: 64'b1010001100111001100100010011100100100101011100011100011100011100;
		8'd220: 64'b0111001001001110101101011110011101110011010101000111000110001110;
		8'd221: 64'b0000001111111001101100110001000011010011111110001101000101001001;
		8'd222: 64'b1000011000100001111111010010010100111100100100010000110110111111;
		8'd223: 64'b0000101110000111001011111100000011001001100100010100001011100000;
		8'd224: 64'b1100111010011100100011101110001011111110111001011010111001101010;
		8'd225: 64'b1010101010101011101000000000110010101100001010011111100010101110;
		8'd226: 64'b0110000101000100010110101100000101111101010000101001001111100110;
		8'd227: 64'b0010011111100000011101110010110101111101001010000010101100101011;
		8'd228: 64'b0100010010001001110001110101111011100100110111101000111100111100;
		8'd229: 64'b0101101100011000010010010101001000110001110111000001100110010110;
		8'd230: 64'b0101111111011100101001110101100000011101110110011110111001010001;
		8'd231: 64'b1000111100011001110001010100001010010011010100011001010010000000;
		8'd232: 64'b0001001110001010110101010110110000000010010110101100010011010111;
		8'd233: 64'b1111111101001010010001111000011001011111001010100111000001111100;
		8'd234: 64'b1111011010010011100010001110000100110100111100111110100100110011;
		8'd235: 64'b0111110100111000011110100001001101110100010100010111011011000100;
		8'd236: 64'b0010001101000011100110101011100000100110000001010100101100111000;
		8'd237: 64'b1010111111010111101011011000001110001011110101101101011000010111;
		8'd238: 64'b1100011011110000001000000101110111100111001111001110110011111000;
		8'd239: 64'b0101011010110011101100001010110110100001001100000000000000111111;
		8'd240: 64'b1110101110100011010101010111110101000010111010000000000111101101;
		8'd241: 64'b1110101101000111111001000001011011111000110011011010010000011100;
		8'd242: 64'b0010101010111000110001111100011110100010110010101010010011001101;
		8'd243: 64'b1111011010010101001010101001100111101000111101110001010010110000;
		8'd244: 64'b0100101101000110000000101111110100100011100001110000101010111010;
		8'd245: 64'b0010000010100101000010011111011010110101111001011011100010001000;
		8'd246: 64'b0100110100001100010000001001110000111100011000110100110111111111;
		8'd247: 64'b1100100100010001010110110010000100000001011110010010100001110101;
		8'd248: 64'b1111010001101101011110100010101001010101101110011011100011001101;
		8'd249: 64'b1110000111010110010001000010000011001010010000100101011010111011;
		8'd250: 64'b0111100100111110111011100001111111011101100010001001010000000101;
		8'd251: 64'b0101100010001111000101100101011010001100110111110111110000010110;
		8'd252: 64'b1011001000110010111010001000010111011010000100100011100010000111;
		8'd253: 64'b1000011000011101110010010101110111010001001001001001100011111110;
		8'd254: 64'b0111101111111001011010101111011010010100111110010011001101111000;
		8'd255: 64'b0000000010000101000101010111100001000001001110010101010101100101;
	endcase;
	return out;
endfunction
function Bit#(256) get_msg_bit_page5(UInt#(4) counter);
	Bit#(256) out = case(counter)
		4'd0: 256'b0010011010000010100001100100110001111001111001100101001010100000101010001111110100100110011100011010101110001001000010110011110010000100000011101011110100101110010000011000010100000111101110011000111000110101100101111000001011011000001001111101010100000100;
		4'd1: 256'b0011111100111101100010010000100111100001010010000001101111010001101110110100101011010000010001010111110010000101101101100101000111000011100111110001011110100011000001010101101111010010101101101100111110000111110110001000001101010110001010011001001011010001;
		4'd2: 256'b1111111100011010111010000000001010100001110011010001010011000001100111011100110101100111001100111010001001010010000010111110101100100110110111001100111101101101010110000101101001000110100110000010101001001111101010100111111011110010000000001110010011110100;
		4'd3: 256'b1011111110101101111111111101001001010010000010110001001110101011110101111000010000101110111011011010000100100011110010001111100101011100100000001110001110001011011110111101000101101000010010000100101101101010011110100011100100010100110101000110000111000101;
		4'd4: 256'b0011100011111011101111110101100111000001010000101001111100101011101000001000111110010000101111010111101101010010111111000110010001110110111100011011111110010011100000010011100101010111001110000111111001001011101010100011101100111111010110100000011011010011;
		4'd5: 256'b0011110011100110101101110010111100101000011000110100110100101010011010001001001101011011101110001101010111101010010001101000011000010010010010011000010101011100001001011010010001101011000001110000100100011110011000101010010111000001011001010110001000011101;
		4'd6: 256'b1101011000110110001010101101001000100100010011100101100101101111001010000110001100001110110000010001101011100010100100100100011111101101000100100000100111011101100010010100000010010101011010000001100011001101110011110100101111001100101110111110001001010111;
		4'd7: 256'b0011010110110101111001010101010011011111100100001001001101100101010111100111100110010100010111100010100110000100110000011001100101000101001101011101010011110000111100000010001101010110011011110010111011101110011010110010111100110110101100000010111011011010;
		4'd8: 256'b0111000010000101110011111101011001010001101110010010000001101111010010001000010101110001101001110011000101001111101011111111000101110010101000011110111111000011010111100011010001011011011011111100111010110101010100111101110110100110111011001100111010111000;
		4'd9: 256'b1011010110111101000000101000110011110110000000000101110010000110001111101100101001010001001111001001010010100000000010111101110010101010011110110010111000000101010010000001000011110010000010110110110100100010001011101011011010010000011100110111111001010101;
		4'd10: 256'b0001001100011010011001001011001010001000110010010100101001101101101001000010111010100000000100011011111011110011010011000111011111010110101010011100101100010101000110101100101111111110000001100111010110110110100101010010111110001110110110011001010100001100;
		4'd11: 256'b0111100101011101010110100010111110101100100001000100111110011010001101100111110101101101110001101011101111110000011111100010010111101110100001001111100000000111110000101001111001011000111101101010010111110000111111100010100000101110101110111000011111101110;
		4'd12: 256'b0011100001011111100111011100110001110100010011011111011101000000101110100001110100010000010010010000110010001010011010011001001001111001110100100101001010001100100111001011011111010101101100101000010111100001001011001110110110100000000100000100000110101000;
		4'd13: 256'b1110111100110111100100000010111110011101111110011100001000001011010100011110000110011110011010101110100100001111110100000100001101111100101001000110010111010010011100000000101111011110010110000010011000010010111110011110101001000010100101010000001111111001;
		4'd14: 256'b0101111001101010010100010110001000111111001110011001101111000001000101111111111000101100101001011111111101000100100001111011011001101000001110110100011010111110110111000111111000011001100111011010010001110110011011110110111111010111111001110011110010010010;
		4'd15: 256'b0011101101101001110100101010001110001000100100000110110110111000101101110000110000111101100110110011101101001001011010111101111101100111111110001110101000110110011111011110011110000101101010010101101101110101111000111011110111000101111101000100111010100100;
	endcase;
	return out;
endfunction
function Bit#(64) get_prev_enc_page5(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1111111111011011111101101101001010111110100110111011111011001000;
		8'd1: 64'b0010111010111110101010011010001011111010111100100010100111000110;
		8'd2: 64'b0011011000000010111011100111010001100011011111110110101100111111;
		8'd3: 64'b1011011011110011000101101001101000111001110111111011001110111001;
		8'd4: 64'b1101000101110011000111111110100011010001111000010111111111101000;
		8'd5: 64'b0101101011111010110110011101011000111000101110101000111011100111;
		8'd6: 64'b0101110011010101101001111110000110111100100011010101010111010001;
		8'd7: 64'b1011011111010100011011100001000000111001100110011101101111010101;
		8'd8: 64'b0101011100100011000010110110100101111111111100010101111100001010;
		8'd9: 64'b0101011110000110101110101000001101000010100011111100100010011100;
		8'd10: 64'b1111100110011000101111001111111010110101001011010011100001001100;
		8'd11: 64'b1001111001110001000111010011010000110001011101111111100110011111;
		8'd12: 64'b1010010001110111110001100101101001000111101101001111011101111010;
		8'd13: 64'b1110110011100110101100011101101000101111110010010011100110011010;
		8'd14: 64'b0101101011010110101010100111001011111110011101110110001011100101;
		8'd15: 64'b0110110100100011011101001010001111110111100101101110010011001011;
		8'd16: 64'b1010010011101111101000111111001111100101101111011101101100010001;
		8'd17: 64'b1110101111100011101001000101001111111000100001100011010001000100;
		8'd18: 64'b1010001110001000111111100110000000111010000010001110011000101000;
		8'd19: 64'b0101111010111111101111111101101011011110110100111011110110100011;
		8'd20: 64'b1010101000011101101011101111101101101011111101111011111111011110;
		8'd21: 64'b0011110111111011111011101011101111101111111110111010111111111111;
		8'd22: 64'b0100100011111010011001100110110001101001011110000011000001101001;
		8'd23: 64'b1011111010011000100001111011110110111101111010010010100110111011;
		8'd24: 64'b1010010110111111110100011011111110001101101101101010100111010111;
		8'd25: 64'b1111111110110101111110111111011110101111011101111110000101110101;
		8'd26: 64'b0001001010011111000001111110110111001111110101111000010010011111;
		8'd27: 64'b0010010111011101010010010010000100100101110010110100111111000111;
		8'd28: 64'b1100101100110010101110100001011110100011111110100000001110000110;
		8'd29: 64'b0110011111101001111101010010111110100001010111011111000111111110;
		8'd30: 64'b0101010010000001001101100100101110010000010001010001110001101001;
		8'd31: 64'b0001101110100110111110111110011101111110101001101101111111101100;
		8'd32: 64'b0100000101111000111000001101100011010001111111100001110111011000;
		8'd33: 64'b1011000101010111011001000110011100100100011101011110101100101110;
		8'd34: 64'b1001010110111010110100110110111100111010101111101110000001101111;
		8'd35: 64'b1011101111111011101011101001110110111000101111111011011110010001;
		8'd36: 64'b1101001101010011101101011111111110011011011010110110111101111111;
		8'd37: 64'b1110011111000011110111111101111011101011110000101011001010010101;
		8'd38: 64'b1100101011001111111111001111111001001101010011001111000011010110;
		8'd39: 64'b1011101111001100111111110001100100110011100010011101101100000001;
		8'd40: 64'b1110110101111110011011101111110011101100110111010100010011111100;
		8'd41: 64'b0011010101010110100111110011001010010100010111001001110000000010;
		8'd42: 64'b1100111101011011011001100001101010000011010100111110010101100111;
		8'd43: 64'b1001101110000101110110011111010010111000101101000101000101011100;
		8'd44: 64'b1111011110011101111101111011110001010111110100110011011111010110;
		8'd45: 64'b0110101111110011110011011001111111000011101110011100011111110011;
		8'd46: 64'b0000110100000100011100111101010100001101001001010100101111100100;
		8'd47: 64'b1110101100011101011011100100100011001000101001100110111011110100;
		8'd48: 64'b1011111110100101011111111001110111111010110010111110111111111101;
		8'd49: 64'b1110101110010011111011100011010011000010100100110100011100110111;
		8'd50: 64'b1000100110001111001000111100111101001101101101011011010101110111;
		8'd51: 64'b1111111010100111101011111001011010111101111000111111110011001111;
		8'd52: 64'b0111010011011110100101010010001110010111000001111100111110010011;
		8'd53: 64'b0101000100010100111101110001110000110000110110000011101011110001;
		8'd54: 64'b1101000111110111110100110101110001111011111111011011011001111001;
		8'd55: 64'b0110011011000111111001001111001010010110111001101100010111110010;
		8'd56: 64'b0100111101000101011111010101000111010101100111000111110011111001;
		8'd57: 64'b0110001101111111011101110110011101100011010111111100111001011100;
		8'd58: 64'b1110001001100011011101110100010011010011010101110110111011001101;
		8'd59: 64'b1010010000111001101111110101001111001110101010010011011111010111;
		8'd60: 64'b1001111110100101001011111010010111001111100001011010011111111101;
		8'd61: 64'b1100110100110101110101000111111011011111111101110111111101100111;
		8'd62: 64'b0110111011000110101001101000000001111010000001101111001101010111;
		8'd63: 64'b1000110010110100011101111011110001111100111110000011111011101110;
		8'd64: 64'b0100010111101111110010000001010100001101111111011101110001111011;
		8'd65: 64'b0111100111011001100110001111100110110011010101011000101010111001;
		8'd66: 64'b0101111110111010010100110111001000111010101010100111010111111111;
		8'd67: 64'b1111111100010111000111110101010101100110010101111111110110010110;
		8'd68: 64'b1001100001100010010111101111110111110111000101101100011011011111;
		8'd69: 64'b1100011101111110000101110111001011100111101101100010101100010010;
		8'd70: 64'b0001110111000100101111000111000110111101110101010100110000101010;
		8'd71: 64'b1011111110111101011110110001011011110111010111100101101110111100;
		8'd72: 64'b1110000100110111011000111001011010000101000100001100001110001110;
		8'd73: 64'b0000110111000101111011000100111100011101010011011011010011000100;
		8'd74: 64'b1111110101111001110001111000001111111111111100011111110101011111;
		8'd75: 64'b0001110011011100010111111110100001000000100111001000100011011111;
		8'd76: 64'b1100110101010110100111111011110111111101110111110001111111111001;
		8'd77: 64'b0110010100011011100010001100111100010100001111010010111111101101;
		8'd78: 64'b1010011111101111100111110111111100010101010010101111110101001011;
		8'd79: 64'b0111100010001111110011111011101001100101101011000000011000111011;
		8'd80: 64'b1111010101110101010111110111110101011100011111011101011111101101;
		8'd81: 64'b1101111010100110101000001100101010111100100011111011010110001001;
		8'd82: 64'b1100100101000000001100000000101011001100111000110111101100101010;
		8'd83: 64'b1010101101100111100111010110010101111011110001110001101111000100;
		8'd84: 64'b1011001010001100100001111110011110110110110001111011111011101100;
		8'd85: 64'b0101011100010001100111110111101100000101110001110011011110010001;
		8'd86: 64'b1011001101100100010011110111011111110110111101101100011101110101;
		8'd87: 64'b1001000011110011100110111001000010010001110110010001011110110101;
		8'd88: 64'b1000111011011111100111010101011110001110101111110000110111001001;
		8'd89: 64'b1011101100100101111000111011111110110111001100111110000101011010;
		8'd90: 64'b1111000011000111111010101100110111111100111111110011011100101111;
		8'd91: 64'b0011100000101110000110000011010100011001001000000001000010010111;
		8'd92: 64'b0000101110111010011011001111101000001111110111101010101011111011;
		8'd93: 64'b0100110110011011011010011111110111101101110110110010101111111010;
		8'd94: 64'b0110101111001101011010010111100001111110100011000100111101101000;
		8'd95: 64'b1101010101110001111100101000110011110000110101011111111000101100;
		8'd96: 64'b0010011110101001111110111110111100101001111111010011111111101100;
		8'd97: 64'b1001111110101010111110101011100010100111001010101111111000000101;
		8'd98: 64'b1110001000010011101001111001101101110011001100100111010000100111;
		8'd99: 64'b0111110111110111011001101101000111010101001101001110010011100100;
		8'd100: 64'b1101111100001001111101011010101111011101001100001101000110111100;
		8'd101: 64'b0011100100100000010001001110011101011001101001100101010110010110;
		8'd102: 64'b0101100011011110011111111111011111111110101111011101111001010111;
		8'd103: 64'b0111011101000011001010111010000011010011011110100110001111010010;
		8'd104: 64'b0110111110001001101100011000111111010011011010111111110111111011;
		8'd105: 64'b0010001001000111011101110000111100001101000101110011110100111011;
		8'd106: 64'b0010111110110011011111101001101110101111011100110010111111011001;
		8'd107: 64'b1011110110110001010001110011100010010001001010000010001001100001;
		8'd108: 64'b1111111100101110011101110110011001011111000011111110111101111111;
		8'd109: 64'b0101101010100110000111111011000011001010111001110100011100100111;
		8'd110: 64'b0110011001101111010001001010110101101100001111010111010011100101;
		8'd111: 64'b0111000110111101101010010111011111111011101011101000101101110000;
		8'd112: 64'b1101000001010011011111100011010010110000110101101111101001110100;
		8'd113: 64'b1001011000001110111111001100100110010011000011000011111110100000;
		8'd114: 64'b1101001000011011001100010010000110011101010111011111011001011011;
		8'd115: 64'b0111100001100101001111111110111101100101111001000010111111101111;
		8'd116: 64'b1000110110101011101111010001100111011101000001011011111100111001;
		8'd117: 64'b0111101100101011101010111010011101001100011001110010100011110011;
		8'd118: 64'b1110110111010010001011001111011001010110110011100010010001000100;
		8'd119: 64'b0101011101110100111100111000001111010111011111001101010001000010;
		8'd120: 64'b0111001111111111010101000110000111100011010111110000010001111111;
		8'd121: 64'b0101101111111111001110100001001111011110011111000001100100111001;
		8'd122: 64'b1011010110010101100110101001101010010011111110111001100101011011;
		8'd123: 64'b0011001001010010001100100000000001101010010100100100101111000010;
		8'd124: 64'b1100101001000100111001111001010011001100011011111010101011101011;
		8'd125: 64'b1011000010111011101000001100110010100000110111101001010010111010;
		8'd126: 64'b0111011001001011001111110001101010110110010001101001011000011010;
		8'd127: 64'b0111101010110111100010111010110100100110101101010101000100100111;
		8'd128: 64'b1100110000111011110111111111010001100110111010111100110111111101;
		8'd129: 64'b0111101111000111111011001110011111101010001011111110011101000110;
		8'd130: 64'b1100000111000111011011111000110110111101100001010101110111100111;
		8'd131: 64'b1000001010110010011001101001100011000110101011111110010110010010;
		8'd132: 64'b1111000110111011010011100110001110000101011011111000111001000110;
		8'd133: 64'b0100001010000011110111001111110101001011110111010111111111011111;
		8'd134: 64'b1011011011111111111001010101110100110010011011110101111111011111;
		8'd135: 64'b1100111000110100111100010101000110111000101001001111110111010010;
		8'd136: 64'b0011011110111001101110111011111111101111000111111010110110111111;
		8'd137: 64'b1001100100111111010010111111100101011001101110101100110100111001;
		8'd138: 64'b0011101100110110001000001100110000111001101011100010100100111100;
		8'd139: 64'b1001111000001110100011001000010110001101001011011010110101010101;
		8'd140: 64'b0111101011101100100101000101101100001010010000101101111011100011;
		8'd141: 64'b1001010010000001010100101110111011010110110001010000111010001100;
		8'd142: 64'b1101111010101000111110111010101010011101101111000010100010101010;
		8'd143: 64'b0110101000111010101000000011001111110011010010100010001001010111;
		8'd144: 64'b0100000110001001011001110110100110100111011110010101101100111100;
		8'd145: 64'b0100101000111001011111110011001100110011001010101111100001110010;
		8'd146: 64'b1010101110111111111101001100101111000001100110111011010001001111;
		8'd147: 64'b0111001001001101010010101111101111010111111111110100011110110111;
		8'd148: 64'b1100001101000010010000100001000001011001011010000000010101011101;
		8'd149: 64'b0010111101101111010111100110011110100111111011101001011011001111;
		8'd150: 64'b1010111010011110101111110110011010111011100010001010111010111110;
		8'd151: 64'b1010101010011111101011101000110110101010000011111100000110001011;
		8'd152: 64'b1111010100111011011011111011101000011101001111001111101001111010;
		8'd153: 64'b1000001010001000010100111010011011110011111111100111110101101010;
		8'd154: 64'b0001101110101010100111111111111110011111101111111001111110101001;
		8'd155: 64'b1101101110110111011101111011010111111011101101010011011110010101;
		8'd156: 64'b1000011010011110100110110010110000101010110110000000110110001110;
		8'd157: 64'b0010101110001010110011101010011110010000001001101110110110000100;
		8'd158: 64'b0011110000010111011001100101111110100010001101101010011000101011;
		8'd159: 64'b1111011110110110110100101001011110010110111101111010011010101010;
		8'd160: 64'b0011101101111110010010010111101101110001111001100111001011111011;
		8'd161: 64'b0101100110101000110101000010110010010111001011110001001000011100;
		8'd162: 64'b1011101110111111011101011100001101111110111101111110101010100111;
		8'd163: 64'b1001000100100101100110010000101111100001101000011010100101001101;
		8'd164: 64'b1111100100100111101100111010010010111110101011000000100110111100;
		8'd165: 64'b0000000000110110011101110010110100011000101011101001000100011111;
		8'd166: 64'b0010001101010111001100110111001110100101111111010011110101010111;
		8'd167: 64'b1101100111000000110101101111011111010110110000011111011011000011;
		8'd168: 64'b0111001011110101001000111111000000100101111001000110111101010011;
		8'd169: 64'b1010010110111010000110111010001000000001111001111100110101111010;
		8'd170: 64'b0110110011101111100000001111111111101111111111101001111010001010;
		8'd171: 64'b0010001110111011111001001010101101110101101010111101011111101011;
		8'd172: 64'b0101011100001010000100001110101101100100010110011001111100101000;
		8'd173: 64'b0011110100000101011010111011011000110011111001110010101011110110;
		8'd174: 64'b1101100111111110001111100101111111111001101101101101111011010011;
		8'd175: 64'b0101001010010000010001111100100001011000101100100101111110101010;
		8'd176: 64'b0100111101010110010110100011011101000010010110100111111010110101;
		8'd177: 64'b0100100001010111101001100100011110001100010010111011110001101001;
		8'd178: 64'b0100011101100011000111110110001011001011011010110101111101111011;
		8'd179: 64'b1011111111011110010110001010110110100000110110100100001000000111;
		8'd180: 64'b0010011011000010101101111001101100101010000101011111111101010101;
		8'd181: 64'b0010000101000101110000010101110110111101011001110110100011010000;
		8'd182: 64'b0100111101111001100001010011101100011011011110010010110110111101;
		8'd183: 64'b0011001111101010011100110100101111101011101010101111111101111010;
		8'd184: 64'b1100101111111101000110111011101011001101111001101011101110000010;
		8'd185: 64'b1001001101111001110101101111110100110111011111111011101110010101;
		8'd186: 64'b0001010101000010011111101111100000000100111001101111010111110100;
		8'd187: 64'b0001011110011000111110011001000110011111010111010011100100111011;
		8'd188: 64'b1011111010101010101010001101101010111111101001101011100110110111;
		8'd189: 64'b1110101101100010001110110110011101110001011001000101101111100100;
		8'd190: 64'b0100001101010011000100000001011101001011000011010100101110010010;
		8'd191: 64'b0101100101101100011001000111111101110011111011000111100101110110;
		8'd192: 64'b0100011101100101000011010110100111111111010000110001100111100000;
		8'd193: 64'b1110011001001011111010011011010011111111100010110111001101110111;
		8'd194: 64'b1110101010000100011101111001110101011111110001001111111011111011;
		8'd195: 64'b1101011110100111010001111111011111000011111100011101011010010110;
		8'd196: 64'b1110111010101100011101101011011100111110001001110010110111110111;
		8'd197: 64'b1111000001001101001010111011110111111000010111111001101100011110;
		8'd198: 64'b0011010001001101101011101011000101110010000011110011100010100000;
		8'd199: 64'b1010001011011011000011001110110110111101100111111100100011011110;
		8'd200: 64'b0001111101110100110101010010110111001000101111011100011100101001;
		8'd201: 64'b1010101110111110001100110010110100111011001111000011001000101011;
		8'd202: 64'b0000001110100101110101011101111111001110100001111011000110000101;
		8'd203: 64'b1010101110101111110110111010111110101000101111110001101111001010;
		8'd204: 64'b1000000110110110101001001111110010101011111101101010011000100110;
		8'd205: 64'b1111011011011000111101110001011011110110110101110100000110011101;
		8'd206: 64'b1110100010101010101011011101110100111011111011001010111011101110;
		8'd207: 64'b0110010101010011111110010111111110010001111100110111101101110111;
		8'd208: 64'b0101001000101010010010100011011011101100010110101101101001000110;
		8'd209: 64'b0110100010101111111000010010100001100000100010101010100110111000;
		8'd210: 64'b0001011111000011010111110110111111110111011001101001110101100000;
		8'd211: 64'b1111010010111100101101010111110110110000010110100110111101001100;
		8'd212: 64'b0000011111100000001111011110100011110111011000010100001001000110;
		8'd213: 64'b1011000100110011011111100111010010110011001101011011101001110100;
		8'd214: 64'b1001111111101010100110110101111110110110011011101110101101111110;
		8'd215: 64'b1110001111001100000010111000001111001101110101111000000110110001;
		8'd216: 64'b0111011000000111111001110000010100000110000010111011111101100110;
		8'd217: 64'b1111001001001010011100000010001001010011010000000111010011000001;
		8'd218: 64'b0010001111011001111110011011011010110001110101001111110111010101;
		8'd219: 64'b1010101101111001100100010011101100100101011100011100011100011101;
		8'd220: 64'b0111011011001110101101011110011101110111010101000111000110001110;
		8'd221: 64'b0000101111111001101100111001000011011011111110001101000101011001;
		8'd222: 64'b1000011000100001111111010010010100111100100100010000110110111111;
		8'd223: 64'b1111101110010111001011111100000011001001110101110100111011100001;
		8'd224: 64'b1100111010111100101011101110001011111110111101011110111001111010;
		8'd225: 64'b1010101010101011101000000010110010101101001010111111100010111110;
		8'd226: 64'b0111000101000100010110111100010101111101010100101001001111100110;
		8'd227: 64'b0010011111101000011101110010110101111101001010000011101100101011;
		8'd228: 64'b1100010010001001110001110101111011100100110111101000111100111100;
		8'd229: 64'b0101101101011000010110010101001001110001110111000001100110010110;
		8'd230: 64'b1101111111011100101011110101101000011101110110011111111011110001;
		8'd231: 64'b1000111110011001110101010100001010011011010100011001111110000001;
		8'd232: 64'b0001011110011010110101010111110100000010010110101101010011010111;
		8'd233: 64'b1111111101001010010001111010011001011111001010100111000001111110;
		8'd234: 64'b1111011010011011100010001110001110110100111100111110100100110011;
		8'd235: 64'b0111110100111000011110100001001101110100010100011111011011000100;
		8'd236: 64'b0010101101000011100110101011101010100110000011011101101100111000;
		8'd237: 64'b1010111111010111101011011000001110001011110101101101011000010111;
		8'd238: 64'b1100111011110000001100000101110111100111001111001111110011111000;
		8'd239: 64'b0111011010110011101100001110111111100001001100000000010000111111;
		8'd240: 64'b1111101111100111111101010111110101000010111011001100000111111101;
		8'd241: 64'b1110111101000111111001000101011011111000110011111110010000011100;
		8'd242: 64'b0011101010111000110001111100011110100010110010111010010011001101;
		8'd243: 64'b1111011011010101001010101011100111101000111101110001010010110001;
		8'd244: 64'b0110101101001110000000101111110100100011100001110010101010111110;
		8'd245: 64'b0010000010100101001010011111011010111101111001011011100011001000;
		8'd246: 64'b0100110100001100010010001101110001111100011000110100110111111111;
		8'd247: 64'b1100100100110101010110110010001100000011011110010010100001110101;
		8'd248: 64'b1111110001101101011110110011101001010101101110011011100011001101;
		8'd249: 64'b1110000111010110110001100010000011001010010000100101011110111011;
		8'd250: 64'b0111101100111110111011100001111111111101100010001101110100101101;
		8'd251: 64'b0101100010001111000101100101011010001110110111110111111001010110;
		8'd252: 64'b1011001000110010111110001000010111011010000100100011100110000111;
		8'd253: 64'b1000011000011101110010010101110111110001011101001001100011111110;
		8'd254: 64'b0111101111111001011010101111011010010100111110010011001101111000;
		8'd255: 64'b0001000010010101000101010111100011000001011110010101010101110101;
	endcase;
	return out;
endfunction
function Bit#(256) get_msg_bit_page6(UInt#(3) counter);
	Bit#(256) out = case(counter)
		3'd0: 256'b0111111001011110011001001110000011010000111000011101011100011000110101010000000110011010110100001101101001110101010111011110110111010001110011110001000011101001100100010110111000100000110101001001100000111110011010110100101010010101101111000111011011101001;
		3'd1: 256'b1110000100111001111101001011011111100000101001000100010011111011010101100100110111010010010110011010011001101000110000111101001010110011010111110010110101100110001110111001111011000110110111011101010010000000100001101110011110111101010110011111110100010001;
		3'd2: 256'b1100000100010000000111101111101101101110011001001111101111100000010101011000100010101000011010100100101110111101101001111110000011111010111001100011110000010011010011001000101001100100111111101011110110100000100111110010000111110110100110111001000010001101;
		3'd3: 256'b1011001100001001010100010110101111000100001000001101110011001000101101001100011110101100011100011000101010011011001010001001011110100111001000101010000100010011001000110011011001010100101100111110010000011100000010111100100100110001001000010100100011010010;
		3'd4: 256'b1011000111000101110111010100111110011010100011000111001111000010100101100000011100110001111001001110101001101111101001010001011101010101001111000011000000100111010110001011101111011111101010010100011001000111110001011010001111000101010111110000000111000000;
		3'd5: 256'b0011110000111010011010101010101000001110111010110000110100111011110100000011011010001111011001010001101000010001101110000111100001010111100110111110001111001111100010111101110111001110111100010000111110000000101011111011111001111101101111010111100011011110;
		3'd6: 256'b1001010110110101111011001100110001101001110110001111000100000000010100001011100110000011100001110000110011001100101000101010001110101001010110110010111111011011101100100100001011000001000010100110010101101010010010001110010000001110011100010111110100010010;
		3'd7: 256'b0100110100011110001010001110100110101100110111010010000000110100111101110100101101110111100110000111111100000011011110010010011001111001010110001010000100011110010011110011111000100111110100110110111110110001010101011100010010000111010101101000100111010000;
	endcase;
	return out;
endfunction
function Bit#(64) get_prev_enc_page6(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1111111111011011111101111101001110111110110110111011111011001000;
		8'd1: 64'b0110111010111110101010011010001011111010111100100010100111100110;
		8'd2: 64'b0011011000100010111011100111111001101011011111110110101100111111;
		8'd3: 64'b1011011011110011001101101001101010111001110111111011001111111101;
		8'd4: 64'b1101001101110011000111111110100111010001111010010111111111101000;
		8'd5: 64'b0101101011111110110110011101011110111010101110101001111111100111;
		8'd6: 64'b0101110111011101101101111110100110111100110011010111010111010101;
		8'd7: 64'b1011111111010101011011111001000111111011100110011101101111010101;
		8'd8: 64'b0101011100111011100110110110101101111111111100010101111100111011;
		8'd9: 64'b0101011110000110101110101000011111000010100011111100101010011100;
		8'd10: 64'b1111110110011000111111001111111110110111001011010011100101101100;
		8'd11: 64'b1001111101110001000111010011011000110101011101111111100110011111;
		8'd12: 64'b1010110101110111111001100111101001100111101101001111011101111010;
		8'd13: 64'b1110111011100110111100011101101000111111110010011011100110111010;
		8'd14: 64'b1101101011010110101010100111011111111110011101111110101011110101;
		8'd15: 64'b0110111100100011111101001010001111110111101101111110010111001011;
		8'd16: 64'b1010011011111111101001111111001111110111111111011101101111010001;
		8'd17: 64'b1110101111100111101001000101011111111010100001100011011001000111;
		8'd18: 64'b1010011110001001111111100110001000111011001010001110011000101000;
		8'd19: 64'b0101111010111111101111111111101111011110111110111011110110101011;
		8'd20: 64'b1010111110011101101111101111101101101111111101111011111111011111;
		8'd21: 64'b1011111111111011111111111111101111101111111110111011111111111111;
		8'd22: 64'b0100100111111010011101100110110001101101011110000011000001101001;
		8'd23: 64'b1011111010011010100011111011110111111111111010011110101110111011;
		8'd24: 64'b1011010111111111110110011011111110001101101101101111100111010111;
		8'd25: 64'b1111111111110111111110111111011110101111111101111110000101110101;
		8'd26: 64'b0001001010011111000001111111111111001111110111111000010010011111;
		8'd27: 64'b0010010111011111011010010010000100100101110011110101111111000111;
		8'd28: 64'b1100101100110010101110100001111110101011111111101000001111100110;
		8'd29: 64'b0111011111101001111101011111111111100001011111011111000111111110;
		8'd30: 64'b0101110010000011001101100100101111110000010001010001110001111001;
		8'd31: 64'b0001101110101110111110111110011101111110101001101101111111111100;
		8'd32: 64'b0101001101111100111100011101100011010011111111111001110111011000;
		8'd33: 64'b1011001101110111011001001110011100100101011101011110101101101110;
		8'd34: 64'b1011010110111110110100110110111100111010101111101111000001111111;
		8'd35: 64'b1011101111111011101111101001110110111100101111111011111110010001;
		8'd36: 64'b1101001101110011111111111111111110011111011110110110111101111111;
		8'd37: 64'b1110111111000011110111111111111011111011110010111111001111010111;
		8'd38: 64'b1100101011101111111111001111111011101111110011101111100111011110;
		8'd39: 64'b1011101111101100111111110001100100110011100010011111111100100001;
		8'd40: 64'b1110110101111110011011101111110011101100110111010100110011111100;
		8'd41: 64'b0011010101011110100111110011001010010100010111001001110000000010;
		8'd42: 64'b1100111101011011111001100101111011000111010100111110010101100111;
		8'd43: 64'b1101101110110101110110011111010110111000101101001101010101011100;
		8'd44: 64'b1111011111011101111101111011111011010111110101110011011111111110;
		8'd45: 64'b1110101111110011110011011001111111000111101110011100111111110111;
		8'd46: 64'b0000110100000100011101111111110100001101001001010100101111101100;
		8'd47: 64'b1110101101011101111011101100110011001100101101100110111011110100;
		8'd48: 64'b1111111111101111011111111101110111111010111011111110111111111111;
		8'd49: 64'b1110101110010011111011100011010111100010110100110110011100110111;
		8'd50: 64'b1000100110001111001000111100111101101101101111011011010101111111;
		8'd51: 64'b1111111010100111101011111001011010111101111011111111110011001111;
		8'd52: 64'b1111010011011110100101010111001111010111000001111100111110010111;
		8'd53: 64'b0101000100010100111101111001110000110000110110000011111011110101;
		8'd54: 64'b1111001111110111111100110101110101111011111111011111011001111001;
		8'd55: 64'b1110011011000111111001001111011010010110111101101100011111110011;
		8'd56: 64'b0100111101010101011111010111000111110101100111000111110111111011;
		8'd57: 64'b0110101101111111011101110110011101100011010111111110111001011100;
		8'd58: 64'b1110001011101111011101110100010011110111011101110110111011001101;
		8'd59: 64'b1010010000111001101111110101011111011110101110011011011111011111;
		8'd60: 64'b1101111110100101011011111011010111001111100001011010011111111101;
		8'd61: 64'b1101110100111101110111010111111111011111111101111111111111110111;
		8'd62: 64'b0111111011000110101101101001001011111010010001101111001101110111;
		8'd63: 64'b1010110011110100011101111011110001111110111110001111111111101110;
		8'd64: 64'b0100010111111111110111000001010100001101111111011101110001111011;
		8'd65: 64'b1111100111111101100110001111100110110111110101111010101010111001;
		8'd66: 64'b0101111110111010011100110111111000111010101010100111010111111111;
		8'd67: 64'b1111111100010111001111110111010101101110011101111111110110010111;
		8'd68: 64'b1011101001100110011111101111110111111111000111101100011111011111;
		8'd69: 64'b1100011101111110110101110111001011101111101101100010101100010010;
		8'd70: 64'b1001111111100100111111000111000110111101110101010101110000101011;
		8'd71: 64'b1011111110111101011110110001011011110111010111100101101110111100;
		8'd72: 64'b1110000100110111111000111001111010000101000100011100011110001110;
		8'd73: 64'b0000110111001101111011001100111110011101110011011111110011000100;
		8'd74: 64'b1111110101111001110011111100101111111111111100011111110101011111;
		8'd75: 64'b0001110011111100010111111111100001000000100111001001100011011111;
		8'd76: 64'b1100110101011110100111111011111111111101110111110001111111111001;
		8'd77: 64'b0110010100011011100010001100111100011100011111010011111111111101;
		8'd78: 64'b1010011111111111100111110111111100010101010010101111110101011011;
		8'd79: 64'b0111100010001111110011111011101101100101101011010101011010111111;
		8'd80: 64'b1111010101110101010111110111110101011100011111011101011111101101;
		8'd81: 64'b1111111010100110101011111101101011111100100011111011010110001001;
		8'd82: 64'b1100100101100000001100000000101011011101111000110111101100101010;
		8'd83: 64'b1110101101100111100111010110010101111011110001110001101111000100;
		8'd84: 64'b1011001010001100100101111110011110110110110001111011111011101111;
		8'd85: 64'b1101011100010101100111110111101100000111110001110011011111010011;
		8'd86: 64'b1011101101110110110011110111011111110111111111101111011101110101;
		8'd87: 64'b1001000011110011110110111001000110011001110110011011011110111101;
		8'd88: 64'b1000111111011111100111011101011110001110101111111000110111001001;
		8'd89: 64'b1111101110110101111100111011111110110111001100111110000101011010;
		8'd90: 64'b1111000111000111111110101101110111111100111111110111011101101111;
		8'd91: 64'b0111100000101110000111000011010100011001011001000001000010110111;
		8'd92: 64'b1110101111111010011011101111101100001111110111101010101111111011;
		8'd93: 64'b0100111110011011011110011111110111101101110111110010101111111111;
		8'd94: 64'b0110101111001101011110011111101001111111111011000100111101101000;
		8'd95: 64'b1101010101110101111100101000111111110001110101011111111001101100;
		8'd96: 64'b0010011111101001111110111110111100111101111111110011111111101101;
		8'd97: 64'b1001111110101010111110101011100010100111101010101111111001100101;
		8'd98: 64'b1110001000010011101011111001101101110011001100100111011000110111;
		8'd99: 64'b0111110111110111011001101101000111010101001101001110010111100100;
		8'd100: 64'b1101111100011001111111011110101111011101001110001101000110111100;
		8'd101: 64'b0011100100100000010001001111011101011011101001110101011110010110;
		8'd102: 64'b0101110011011111111111111111111111111110111111111101111001010111;
		8'd103: 64'b0111011101000011001010111010001011110011011110100110001111010110;
		8'd104: 64'b1110111110001011101100011000111111010011011010111111110111111011;
		8'd105: 64'b0010011011000111011101110010111100101111001101110111110100111011;
		8'd106: 64'b1010111110111011011111101011111110101111011100110010111111011001;
		8'd107: 64'b1011110110111001010011110111100010010011001110010010011001100001;
		8'd108: 64'b1111111100101111011101110110011011011111010011111111111101111111;
		8'd109: 64'b0101101010100110000111111111011011001010111001110110011100110111;
		8'd110: 64'b0110011001111111010001011010110101101101001111010111011011100101;
		8'd111: 64'b0111001110111101111010010111011111111011101011101100111101110110;
		8'd112: 64'b1101100001010111111111100011010010110100110101111111111011110101;
		8'd113: 64'b1001011000001110111111001110100110110011000011001011111110101000;
		8'd114: 64'b1101001000011011001100110010000110011101010111011111011001111011;
		8'd115: 64'b0111100111100101011111111110111101110111111001000010111111111111;
		8'd116: 64'b1011111110101011101111010011100111011101000001011011111100111001;
		8'd117: 64'b0111101100101011101010111110111101001100111001111010111011110111;
		8'd118: 64'b1110111111010111001011001111011001010111110011100010111001000100;
		8'd119: 64'b0111011101111101111100111000001111010111011111001101010101000011;
		8'd120: 64'b0111001111111111110101010111001111100111011111110000011001111111;
		8'd121: 64'b0101101111111111001110100001001111011110011111000001100100111101;
		8'd122: 64'b1011010110011101100110101001101010010011111110111001101101011011;
		8'd123: 64'b0011001001010010001100100000000101101111010101100110101111001010;
		8'd124: 64'b1100101001001100111001111001010011001100011011111010101011101011;
		8'd125: 64'b1011010010111011101010001100110010100100110111101001010110111011;
		8'd126: 64'b0111011001001011001111110001101010110111010001111011011010011010;
		8'd127: 64'b0111111110110111100010111010110100100110111101010101000101100111;
		8'd128: 64'b1100110001111111110111111111010011101111111011111110111111111111;
		8'd129: 64'b1111101111001111111011101110111111111010111011111110011101011110;
		8'd130: 64'b1101000111000111011011111000110111111101100011110101111111100111;
		8'd131: 64'b1100001010110010011001101101100011010111111011111110111110010010;
		8'd132: 64'b1111000110111011110011100110011111000111011111111000111001100110;
		8'd133: 64'b0100001010000111111111001111110101001011110111110111111111011111;
		8'd134: 64'b1011011011111111111101010101110101110011011011110101111111011111;
		8'd135: 64'b1100111010110100111100111101100110111010101011001111110111010010;
		8'd136: 64'b0011111110111101101111111011111111101111000111111011110111111111;
		8'd137: 64'b1001100100111111010010111111110101011001101110101100110100111011;
		8'd138: 64'b0011101100110110001010001101110000111001101011100010100100111100;
		8'd139: 64'b1001111000001110100111101000010110011101011011011110111101111101;
		8'd140: 64'b0111101011101110100101000101101100101010010100101101111011110111;
		8'd141: 64'b1001010011000001010100111110111011110110110001010000111010001100;
		8'd142: 64'b1101111010101110111111111010101010011111101111000011100010101010;
		8'd143: 64'b0111101000111010101101000011001111110011010010100010001001010111;
		8'd144: 64'b0100100110001001011001110110100110100111011110010101101100111110;
		8'd145: 64'b0101101000111011111111111011001100110011001110101111100101110011;
		8'd146: 64'b1011101111111111111101001101101111000001100110111011011001001111;
		8'd147: 64'b0111011101101111010110101111111111110111111111110100111110111111;
		8'd148: 64'b1100001101101010010000111011000001011001011010000000010101011111;
		8'd149: 64'b1110111101101111010111100110011111100111111011101101011011001111;
		8'd150: 64'b1010111010011110101111111110111010111011111010001010111011111110;
		8'd151: 64'b1010111010011111101011101000110110101010100011111110100110001011;
		8'd152: 64'b1111010101111011011011111011101000111101001111111111101101111010;
		8'd153: 64'b1011001011001000010100111010011011110011111111100111111101101010;
		8'd154: 64'b0101111111101110100111111111111110011111101111111001111110111101;
		8'd155: 64'b1101101110110111111101111011110111111011101101010011011110110101;
		8'd156: 64'b1010111010011110100110111110110100101010110110000000110111001110;
		8'd157: 64'b0010101110001011110011101010011110010000001001111110110110000100;
		8'd158: 64'b0111111000011111011001110111111110100010001101101010011000101111;
		8'd159: 64'b1111011110110111110101101001011110110110111101111010011010101011;
		8'd160: 64'b0111101101111110111010111111111101111101111101101111001011111011;
		8'd161: 64'b0111100110111000111101100010110011011111101011111001001100011100;
		8'd162: 64'b1111101111111111011101011100011101111111111101111110101010100111;
		8'd163: 64'b1001000101110101101110011000101111101001101010011110100101001101;
		8'd164: 64'b1111101110101111101100111010110010111111101011000010100111111100;
		8'd165: 64'b0000010000110110011101110010111100011000101011101001001110011111;
		8'd166: 64'b1011001101010111001100110111001110100101111111110011110101010111;
		8'd167: 64'b1101101111100011111101101111011111010111110000011111011011000111;
		8'd168: 64'b0111001011110111101001111111000010100101111101000110111111010011;
		8'd169: 64'b1010110110111011000110111011001000000011111001111100111111111010;
		8'd170: 64'b0111110011101111100000001111111111101111111111111001111110011010;
		8'd171: 64'b0110001110111011111001001010101101110101101010111101011111101011;
		8'd172: 64'b0111111100001010000100001110101101100100010110011001111100101000;
		8'd173: 64'b0011110100110101011010111011011000110111111001110010101011110110;
		8'd174: 64'b1101100111111110001111101101111111111001101101101101111011010011;
		8'd175: 64'b0101011010010000010001111100100001011000101100100111111111101010;
		8'd176: 64'b1100111101010110010110100011011101001010010110100111111010110101;
		8'd177: 64'b1100100001010111101001100100011110001100010010111011110001101001;
		8'd178: 64'b0110011101101011000111110110001011011011011010110101111111111011;
		8'd179: 64'b1011111111011110110110001010110110101010110110100100101000000111;
		8'd180: 64'b0010111011100110111111111101111100101011100101011111111101010101;
		8'd181: 64'b0010010101100111110011010101110110111101011001110110101011010000;
		8'd182: 64'b1110111101111001101011010011101100011111011110010010110110111101;
		8'd183: 64'b0011001111101111011101111100111111101111101010101111111101111010;
		8'd184: 64'b1100101111111111000110111011101011011101111011101011101111000011;
		8'd185: 64'b1101001101111001111101111111110110110111011111111111101110110101;
		8'd186: 64'b0001010101000110011111101111100000110101111001101111010111110100;
		8'd187: 64'b0001011110011000111110011011101110111111011111010011100110111011;
		8'd188: 64'b1011111010111110101010001111111110111111101001101011101110111111;
		8'd189: 64'b1111111101100010001110110110011101110001011001101101101111110110;
		8'd190: 64'b0100101111010011000101000011011101001011000111110100101111010010;
		8'd191: 64'b0101100101101100011101000111111101110011111011000111100101110110;
		8'd192: 64'b1100111101100111000011011110100111111111010100110011101111100001;
		8'd193: 64'b1110011001001011111111011011010011111111100010110111001101110111;
		8'd194: 64'b1110111110001101011101111001110111011111110011011111111011111011;
		8'd195: 64'b1111011111110111110001111111011111010111111100011101011010011111;
		8'd196: 64'b1110111010101111011111101011011100111110001001110010110111110111;
		8'd197: 64'b1111100001001101111010111011111111111100011111111011101100111110;
		8'd198: 64'b0111010001101101101011101011000101110010100011110011101010100001;
		8'd199: 64'b1010101111111011001011001110110110111101100111111100100011011110;
		8'd200: 64'b0101111101111100110101010111110111001100101111011101011101101001;
		8'd201: 64'b1010101110111110001100110010111110111011001111000011001000101011;
		8'd202: 64'b1000001110110111111101111111111111011110100001111011010110000101;
		8'd203: 64'b1011111110101111111110111110111110101001101111110001101111001010;
		8'd204: 64'b1010000110111111111001001111110011101011111101101010011100101110;
		8'd205: 64'b1111011011011000111101110001011111110110110101110100001110011101;
		8'd206: 64'b1111100010101110101011011101110100111011111011001010111011111110;
		8'd207: 64'b0111111101010111111110110111111110010101111110111111101101111111;
		8'd208: 64'b0111011010101010010010100011011111101110011110101111101001000110;
		8'd209: 64'b0110110010101111111000010010100001100000101011101010110110111100;
		8'd210: 64'b0111011111100011010111110110111111110111011001111001110101101000;
		8'd211: 64'b1111010010111110101101011111110110110000010111100111111101001100;
		8'd212: 64'b0000011111100000011111011110100011110111011000010100001011000110;
		8'd213: 64'b1011100100110011111111110111010010110011011101011011111001110100;
		8'd214: 64'b1101111111101011101111110101111110110110011011101111101101111111;
		8'd215: 64'b1110001111001100100010111011001111011101110101111000000110110001;
		8'd216: 64'b0111011001000111111001110000010100000110010010111011111101100110;
		8'd217: 64'b1111111001001010011100100010101001010011010001100111010011000011;
		8'd218: 64'b0111101111011101111110011011111010110001110101011111110111010101;
		8'd219: 64'b1010111101111101110101010111101100100101011100011100011100011101;
		8'd220: 64'b0111011011001110101101011110011101110111010101010111000110001111;
		8'd221: 64'b0001101111111001111101111101100111011111111110011101000101111111;
		8'd222: 64'b1001111000100001111111010010110100111100100100010000110110111111;
		8'd223: 64'b1111101111010111101011111100000111001001110101110100111111101001;
		8'd224: 64'b1101111011111100101011101110001011111110111111011110111001111110;
		8'd225: 64'b1010101010101011101000000010111011101111001010111111100010111110;
		8'd226: 64'b0111010101000100010110111100010101111111011101101001001111100110;
		8'd227: 64'b0010011111101001011111110011111101111101001010001011101100101111;
		8'd228: 64'b1100010010101101110101111101111111100110110111101001111100111100;
		8'd229: 64'b0101101101011000010110011101001101110011111111000001110111010110;
		8'd230: 64'b1101111111011100101011110101101000011101110110011111111011110001;
		8'd231: 64'b1001111110111001110101110100001110011011010100011001111110000001;
		8'd232: 64'b0001011110011010110101110111110100000010010111101101010011010111;
		8'd233: 64'b1111111101001010010001111010111001011111001010100111000001111110;
		8'd234: 64'b1111011011111011101011001110001111111100111110111110100100110111;
		8'd235: 64'b0111110100111000011110100101001101111100010100011111011011000100;
		8'd236: 64'b0010101111000011100110101011101010100110000011111101101100111000;
		8'd237: 64'b1010111111010111101011111000001110001011110101101101011111010111;
		8'd238: 64'b1101111011111000011100000101110111100111111111001111110011111100;
		8'd239: 64'b0111011010110011101100011111111111100001001100011000010000111111;
		8'd240: 64'b1111111111101111111101010111110111111010111011001110000111111101;
		8'd241: 64'b1111111111000111111001100101011111111010110011111110110000111100;
		8'd242: 64'b0011101110111010110001111100111110100110110010111010010111001111;
		8'd243: 64'b1111111011110101001011101011100111101100111101111101010110110001;
		8'd244: 64'b0110101111001110000000101111110100101111110011110010101010111110;
		8'd245: 64'b0010000010100111001010011111011010111101111001011111100111001100;
		8'd246: 64'b0100110101001100110011011111110001111100011110110100110111111111;
		8'd247: 64'b1100100101110101010110110011101100010011011110010010101001110101;
		8'd248: 64'b1111110001101101011111110111111011010101101111011011101111011101;
		8'd249: 64'b1110000111010110110001100010000011001010010101100101011110111111;
		8'd250: 64'b0111111100111110111111100001111111111101100111001101110100101101;
		8'd251: 64'b0101100110011111010101100101011011001110110111110111111001010110;
		8'd252: 64'b1011101001110010111110011000010111011010001100100011100110010111;
		8'd253: 64'b1001011000011101110010011101110111110001011111101001100011111110;
		8'd254: 64'b0111111111111011011110101111011110010110111110010111101101111000;
		8'd255: 64'b0101000011010101000101010111110111110001011110011101010101110101;
	endcase;
	return out;
endfunction
