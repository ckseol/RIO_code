function Bit#(64) get_output(UInt#(8) counter, UInt#(3) page_num);
	Bit#(64) enc_output = case (page_num)
		3'd0: get_output_page0(counter);
		3'd1: get_output_page1(counter);
		3'd2: get_output_page2(counter);
		3'd3: get_output_page3(counter);
		3'd4: get_output_page4(counter);
		3'd5: get_output_page5(counter);
		3'd6: get_output_page6(counter);
	endcase;
	return enc_output;
endfunction

function Bit#(64) get_output_page0(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b0000110010000000000000000000000000010100100100000000100001000000;
		8'd1: 64'b0010000000000000000000000000000000111000010000100000100001000000;
		8'd2: 64'b0000000000000000010000000110000000000000011000000010100000000000;
		8'd3: 64'b0000001000000010000001000000000000001000100010000010000100100000;
		8'd4: 64'b0101000000000000000001010000000010000000000000000000000011000000;
		8'd5: 64'b0000001000110000000000001100011000000000101000100000000000100001;
		8'd6: 64'b0001010010010100000000000000000000000000000000000000000000000000;
		8'd7: 64'b0000000000000100000001000001000000000000000010000100000101000000;
		8'd8: 64'b0100000000100011000000100000000000000100000100000001001000000000;
		8'd9: 64'b0100011000000000000000001000000000000000000000101000000000000000;
		8'd10: 64'b0011000100010000101000001001000000000100000000000000000000001000;
		8'd11: 64'b1000000001000001000000000000000000000000000000000010100000000001;
		8'd12: 64'b0000010000000000000000000000000000000001000100000010000000000010;
		8'd13: 64'b0000000000000000000000000000101000000001110000010010000000000010;
		8'd14: 64'b0100100000000000100000000000000010000000000000110000001000000101;
		8'd15: 64'b0010000000000001000101000000000010000000000000000010000010000000;
		8'd16: 64'b0000000011000000000000000000000011100000101100000000000000000001;
		8'd17: 64'b0000100000000000000000000001000100001000000001000001000001000000;
		8'd18: 64'b1000000010000000001000100000000000000000000000000000011000100000;
		8'd19: 64'b0100101000010001000010100000000010001000100000000000000000000000;
		8'd20: 64'b0000000000000000000000100000100100000000000000010000001001010010;
		8'd21: 64'b0000000111000000100000000011000100000011000000000000100000100101;
		8'd22: 64'b0000000000000000000001000000100000001000000010000000000000000000;
		8'd23: 64'b0000110000000000000000000000000000010000000000010000000000100000;
		8'd24: 64'b1000000000110010100000000000000000000100000000000000000110000001;
		8'd25: 64'b1000001000000000010000100000000100001010000000000000000000000000;
		8'd26: 64'b0000000010000101000000010000000000000011000000010000010000000001;
		8'd27: 64'b0000010010000100000000010000000000000000000000100000000100000010;
		8'd28: 64'b0000000000000010000100000000000100000001000000000000001000000000;
		8'd29: 64'b0110000010000000000100000000000000000000010000000001000000000000;
		8'd30: 64'b0000000000000000000000100000000000000000000001010000000000100000;
		8'd31: 64'b0000000100000010000000001110000000001000000001100000000000000000;
		8'd32: 64'b0000000001010000011000000000100000000000000100000000000000000000;
		8'd33: 64'b0000000000010101001000000000001000000000010000001100000000000000;
		8'd34: 64'b0000000100100000010000000100000100010000000101000000000000100001;
		8'd35: 64'b0000000100010000000000000000100000000000000000001000001010000000;
		8'd36: 64'b0000001000000000100101010000001000001000010000000000001000000000;
		8'd37: 64'b0110000010000001000000000000000000000000110000000001000000000100;
		8'd38: 64'b1000000001000000000000000000001000000000000001000000000000010100;
		8'd39: 64'b0000000010000000000010000001000000000000100000001100000000000000;
		8'd40: 64'b0100000000000000000000000001000000100000010001010000010001000000;
		8'd41: 64'b0000000100010000000000110000000000000000000010000001000000000000;
		8'd42: 64'b0000000000000000000000000000100000000000000000000100000000100000;
		8'd43: 64'b1001000110000000000000000000010000000000000000000001000001000000;
		8'd44: 64'b0101010000000001001100100000100000000010100100010000000000010000;
		8'd45: 64'b0000100000000000110000001000000000000010000000000000000010010010;
		8'd46: 64'b0000000000000000000000000000000100000100000000000100001111000000;
		8'd47: 64'b0100100000000000000010000000000000000000001000000000000010010000;
		8'd48: 64'b0000000000100000000000010000000001110000000000001000000001001000;
		8'd49: 64'b1000000000000001001000000000000000000000100100010000011000000000;
		8'd50: 64'b0000000000001111000000000000010100001000000001000000000000000000;
		8'd51: 64'b1000111000000010000010000000000000000000000000001010000000000000;
		8'd52: 64'b0100010000000000000000000000000000000010000001001000000000010000;
		8'd53: 64'b0100000000010100010000010000000000000000000000000000000000000000;
		8'd54: 64'b0100000000000000000000010000000000100000100001001000000001100000;
		8'd55: 64'b0000000000000010110000001100000000000000000000000000010000000000;
		8'd56: 64'b0000000100000001000000000000000001010000000000000101010000000001;
		8'd57: 64'b0100001000000000000000010010000100000010000000010100010001000000;
		8'd58: 64'b1000000001000000000000000000000000000010000001010010001000001101;
		8'd59: 64'b0000000000101000000010100000000000000000000000000001000101000000;
		8'd60: 64'b0000000100000000001000001010000011000000000000000010000000000000;
		8'd61: 64'b0000100000000000000100000101000000001010111000000101101000100000;
		8'd62: 64'b0000010000000010000000001000000001000010000000000100001000000000;
		8'd63: 64'b0000000000010000001000000010000000001000000000000001000000000000;
		8'd64: 64'b0100000101000000100010000001000000001000100000001000010000000000;
		8'd65: 64'b0000000100011000000000001001000000000000000100000000000000000000;
		8'd66: 64'b0000000000000010000000000000000000010000000000000011000100000000;
		8'd67: 64'b0000000100010000000001100000000000000100000000001010000010000100;
		8'd68: 64'b0000000001000000010000100010000000000000000100000000000001001000;
		8'd69: 64'b1000010000000100000000000000000000000100000101100000000000000000;
		8'd70: 64'b0000000000000000000101000000000000010000010000000100100000001000;
		8'd71: 64'b0010000110000100010110000000001000010010000000000000001000000100;
		8'd72: 64'b1000000000000111010000000000010000000000000100000000000000000000;
		8'd73: 64'b0000000000000000000001000000111000000100000000000000000011000000;
		8'd74: 64'b0011100000000000000000100000000100000010000000001000000000000000;
		8'd75: 64'b0001000010000000000000010000000000000000100001001000000000011000;
		8'd76: 64'b0000000000000000000000010001000100000101000010110001000000000000;
		8'd77: 64'b0000000000000000100010000100000000010000000100000000001000001000;
		8'd78: 64'b0000000000001010000000010100010100000000000010100110000000000000;
		8'd79: 64'b0000000000000100000000001000100001100000000011000000000000000000;
		8'd80: 64'b0000010000000000000000010000010001001000000100011000000001000100;
		8'd81: 64'b0001000010000000000000000000001000011000000000000000000000000000;
		8'd82: 64'b0000000000000000001000000000001000001000000000100000100000100000;
		8'd83: 64'b0000000000000001100001000100000100100000000000010000000100000000;
		8'd84: 64'b0000001000001000100000000100000000000000000000010001011000001000;
		8'd85: 64'b0000001000010001000000000000000000000100100001000000000000000000;
		8'd86: 64'b0010000101000000000011010000000010000010010000000000000100000000;
		8'd87: 64'b0001000010010000000000000000000000000000000010000000010000100100;
		8'd88: 64'b0000001010000010000010010000011000000000000000000000010100000000;
		8'd89: 64'b0001000000000000001000000000001000000000000000000000000100001000;
		8'd90: 64'b0100000000000100000010000000000010110000000000100000001000000000;
		8'd91: 64'b0000000000000000000000000000010000010000000000000001000000000001;
		8'd92: 64'b0000100000100000000000000000100000000010110010100010000000010010;
		8'd93: 64'b0000000100000011010000000001100000000000000100000000000000100010;
		8'd94: 64'b0000000000000000000010000000000000100000000000000000001100000000;
		8'd95: 64'b1000000000100000001100000000010000100000000000000000000000000000;
		8'd96: 64'b0000000010000000000000010010000000000000000000000000000000000000;
		8'd97: 64'b0000000000001000001000001000000000000000001010000010000000000001;
		8'd98: 64'b0000000000000000100000100001000100100000000000100100010000000000;
		8'd99: 64'b0000000010000100000000000100000100000000000000001010010000000000;
		8'd100: 64'b0000100000000001100000011000100100000000000000000000000010100000;
		8'd101: 64'b0011000100100000000000000010000001010000000001000100000000000000;
		8'd102: 64'b0000000000000100010000100000010000001000000000001000100000000010;
		8'd103: 64'b0001010000000000000000000010000000000010001000100100001000000010;
		8'd104: 64'b0000001000000000000100000000000000010000010000011111000001001001;
		8'd105: 64'b0010000000000000000000000000001000000000000000010000000000000000;
		8'd106: 64'b0000010000110000000000000001000000000100001100010000000010000001;
		8'd107: 64'b0000000010100001000001000001000010000001000000000000000000000000;
		8'd108: 64'b1000010000000000000100100000001000000000000000000000100100001000;
		8'd109: 64'b0000000010000100000010000000000000000000001000010000001100000011;
		8'd110: 64'b0000001000000010010000000000000001100000000110010001000000100000;
		8'd111: 64'b0001000000000000000000010000000001101000000010001000000000000000;
		8'd112: 64'b0101000000000000000100000001000000000000000001001000001000000000;
		8'd113: 64'b1001000000001000000000001000000000000010000001000000000100000000;
		8'd114: 64'b0100001000000000001100000010000000000000000000001001000000000010;
		8'd115: 64'b0010100000000000000001010000100100000001000000000000000000001011;
		8'd116: 64'b0000000000001000001101000001000110001000000000000001000100000000;
		8'd117: 64'b0000000100000011001000000010010100000100011001000000000001000010;
		8'd118: 64'b1010000000000000000001000100000000000000000000000010000000000000;
		8'd119: 64'b0000011000100000000000010000001100000001001001001000000000000000;
		8'd120: 64'b0010000010010001010101000000000011000000000000000000010000000000;
		8'd121: 64'b0000000001010000001010000000000101001000000000000000100100010000;
		8'd122: 64'b0000000000000000000000000000000000000000001110010001000000000000;
		8'd123: 64'b0000001000000000000000000000000000000000000000100000000000000000;
		8'd124: 64'b1000000001000000001000000001000000000100000001100000001010001001;
		8'd125: 64'b0000000000010010000000000000010010000000000000000000000000100000;
		8'd126: 64'b0000000000000001000000010000000000010010000001100000010000000000;
		8'd127: 64'b0100000000000000000000000000000000000000001100010000000000100000;
		8'd128: 64'b0000000000110000000111000000000001100100100000001100000100100101;
		8'd129: 64'b0000000110000000001000001000010100000000000001000010000001000000;
		8'd130: 64'b0000000000000001000010000000100000000001000001000001000000100000;
		8'd131: 64'b1000000000100000000000000000000010000000000000100100000000000000;
		8'd132: 64'b0000000010000000000000000110000010000000000000010000000000000010;
		8'd133: 64'b0100000010000000000000000000110000001000000000000000000000000100;
		8'd134: 64'b0011000000101001000001010000000000010000000000100000000001000100;
		8'd135: 64'b0100000000000000000000000100000000000000001000001000010010010000;
		8'd136: 64'b0000000100010000000000010000110010001000000000000000000000010100;
		8'd137: 64'b0000100100100010000000001001000000010000100010000000100000010000;
		8'd138: 64'b0010001100000100000000000100000000000001000000100000000000000000;
		8'd139: 64'b1000000000000100000001001000000010000001000000000010000101000000;
		8'd140: 64'b0011000000000000100100000000000000000000000000001000000000100000;
		8'd141: 64'b0001010010000000010000100010010010000000010000000000000010000000;
		8'd142: 64'b0000010010001000000000010010100000000000000000000000000000100000;
		8'd143: 64'b0000100000000000000000000010000110000010000000000000000000010100;
		8'd144: 64'b0000000010000000010000000000000010100001000000000000000000000100;
		8'd145: 64'b0000000000000000010001100000000100010001001000000000000000010000;
		8'd146: 64'b0000001000100000000001000000000000000000000000000010000000000000;
		8'd147: 64'b0000000000000000010000000010000001000010100000000000000000000101;
		8'd148: 64'b0000001001000010000000100000000000000001001010000000000000000000;
		8'd149: 64'b0000000000001000000000000100000010100000010010100000000001000000;
		8'd150: 64'b0010100000000100001000010010000010001011000000000000011000000000;
		8'd151: 64'b0010000000000100100000000000100100000000000000101100000000000000;
		8'd152: 64'b1010000000110001000000010000000000000000001000000000000000000000;
		8'd153: 64'b0000001000000000010000000010000000000000100000100000000100000010;
		8'd154: 64'b0000000000000000000101010100000000000010100000000001001000000000;
		8'd155: 64'b0000000010110000000000010000010000010001000000000001001100010000;
		8'd156: 64'b0000000000010000000000000000100000000000100000000000000000000100;
		8'd157: 64'b0010000100000000000000000000000000000000000000000000010010000100;
		8'd158: 64'b0000100000000010000000000000000000100000000101000000001000001010;
		8'd159: 64'b0010000010000110000100000000000010010000101100001000011000001000;
		8'd160: 64'b0000000000000000000000000011000000100000000000000010000000100010;
		8'd161: 64'b0000000000100000000000000000100000000000001000000000000000010000;
		8'd162: 64'b0000000010000000000000000000000000010000100000110000000010000010;
		8'd163: 64'b0000000100000100000000000000100000000000000000000000000100000000;
		8'd164: 64'b0000000000000000000000000000010000000100001001000000000110111100;
		8'd165: 64'b0000000000000000010100010000010100000000101000100000000000010000;
		8'd166: 64'b0000000000000100001000000000000010100001100000010001000000010010;
		8'd167: 64'b1000100000000000000000000000001011000000000000010010010001000000;
		8'd168: 64'b0000000000000001000000100010000000000000000000000000100101000000;
		8'd169: 64'b0010010010100000000000000000000000000000011000000100000000000000;
		8'd170: 64'b0000100000000000000000000011010110000010011000001000110010001000;
		8'd171: 64'b0010000000001000000000000010001100000100100000110001000001001000;
		8'd172: 64'b0000001000000000000000000000100000000000000000000000000000000000;
		8'd173: 64'b0000000000000100011000000000010000000000011000000000001000000000;
		8'd174: 64'b0001000000000000000010100000000100000001101000000001000000010000;
		8'd175: 64'b0100000000010000000000101000000000000000000000000001000000000000;
		8'd176: 64'b0000000000000100000010000000000000000000000000000010010000100001;
		8'd177: 64'b0000000000010100000000100000000010000000000000000000000001001000;
		8'd178: 64'b0100010000100000000100000000000000001000001010100000000000010001;
		8'd179: 64'b0000000100000010000100001000100100000000100010000000000000000000;
		8'd180: 64'b0000000010000000100100010000000000001010000000000000001000010000;
		8'd181: 64'b0010000001000000000000000000000000100000010000000100000000010000;
		8'd182: 64'b0100000100000001000000000000000000000010000010000010000000000001;
		8'd183: 64'b0000001001000000000000010000001000000000101000001000000101001000;
		8'd184: 64'b0000000001001001000010001011100001000000000001000000001000000000;
		8'd185: 64'b0000001101000000010100000001010000000100000000000000001000000000;
		8'd186: 64'b0000000000000010000001000100100000000000000000000000010000000000;
		8'd187: 64'b0000011100000000110100010000000000000000010000000000000000100000;
		8'd188: 64'b1001000000001000100000000001000000000000000000100010100100000101;
		8'd189: 64'b1010000000000000000000000000000000000000010000000000001010000100;
		8'd190: 64'b0000000000000001000000000001000000000001000010000000000000000000;
		8'd191: 64'b0001000000000000001000000100000000100000010000000000100101000000;
		8'd192: 64'b0000000000000000000000010110000010000000010000000000000001000000;
		8'd193: 64'b1100000001001000001000000000000000000100000000010000001000010000;
		8'd194: 64'b0100000000000000000101010000000000000000100001000000000000100000;
		8'd195: 64'b0100001110100000010000000000001011000010001000000000000000000000;
		8'd196: 64'b0000011000000000000101000000000000001000000000000010000100010100;
		8'd197: 64'b0010000000001101000000100001000001000000010000000001100100001000;
		8'd198: 64'b0000000000000000000001100001000000000000000010010000000000000000;
		8'd199: 64'b0000000001000001000000000000000010000000100000000100000010001000;
		8'd200: 64'b0001010000100100000000000000110100001000000100000000000000001000;
		8'd201: 64'b0000001100100000000000000000010000110000000001000000001000001000;
		8'd202: 64'b0000000000000100100000011000010000000000000000100000000000000000;
		8'd203: 64'b0000000000100000010000010000000000001000000000010000000001000000;
		8'd204: 64'b0000000100000000000001000010000000100001000000100010000000100010;
		8'd205: 64'b0001000000000000000000000000000010100000000000000000000100000100;
		8'd206: 64'b1000000000000000001001000000100000000000000000000000100000000010;
		8'd207: 64'b0010000000000001000100000010011010000000000100000001000101000011;
		8'd208: 64'b0100000000000000010000100000000000000000000000000100000000000000;
		8'd209: 64'b0000100000000100000000010000100000000000000010001010100010000000;
		8'd210: 64'b0000000000000000000010000000000101100000001000000000010000100000;
		8'd211: 64'b0010000000000000000000010100000000010000000000000010100000000100;
		8'd212: 64'b0000010100000000000000000010000001010100000000000000000001000000;
		8'd213: 64'b0001000000000000001000000000000000100010000000001000100001010000;
		8'd214: 64'b0001000010000000100000000000000000000110000000001000001000001000;
		8'd215: 64'b1000001001000000000000100000000000000000100000101000000110000000;
		8'd216: 64'b0000000000000000100001000000000000000010000000010001000000000000;
		8'd217: 64'b0101000001000000000000000000000000000000000000000001000000000001;
		8'd218: 64'b0010001000011000000000001010000000000000100000000000100001010000;
		8'd219: 64'b0010000000000000000000010000000000100000000100000100000000000000;
		8'd220: 64'b0000000000000000001000001000010000010000010000000000000100000100;
		8'd221: 64'b0000000010000000000100000000000010010010001000000000000000000000;
		8'd222: 64'b0000001000000000001100000000000100100000000000000000000000010110;
		8'd223: 64'b0000000010000100000000010000000000000001000100000100000000000000;
		8'd224: 64'b1000001000010000000000000010001011000000110000010000110000000010;
		8'd225: 64'b0000000000001000100000000000010010000100000000000001000000100000;
		8'd226: 64'b0000000000000000000000000000000001100001010000000001000010000000;
		8'd227: 64'b0000000000100000000000000000000000000100000000000000100000000001;
		8'd228: 64'b0000000000000000010000000101100000000100010001001000000000011100;
		8'd229: 64'b0000000000010000000010000001000000000000000000000001000100000000;
		8'd230: 64'b0000000000000100000000000000100000000001000000001010001001000000;
		8'd231: 64'b0000011000000000000001010000000000000000000000010000000000000000;
		8'd232: 64'b0000001010000000100000000000000000000000000000100000000000000100;
		8'd233: 64'b0010000000000010000000000000000000010101000000000100000000011100;
		8'd234: 64'b0000001000000001000000000010000000100100000000110000000100000000;
		8'd235: 64'b0100000100000000000100000000001000000000000000000000001010000000;
		8'd236: 64'b0000000000000000000100000000100000100000000000000000000100000000;
		8'd237: 64'b1000000000000000000000000000001000001000010001100000000000000000;
		8'd238: 64'b0100010000000000001000000001000000100111000010000000000000001000;
		8'd239: 64'b0000000010110000000100000000000100000000000000000000000000001001;
		8'd240: 64'b0000001000000000000000000101000100000000101000000000000000101001;
		8'd241: 64'b0000000000000000000000000000001000001000110001000000000000000000;
		8'd242: 64'b0000000000010000010001101000010100100000000010000000000000000001;
		8'd243: 64'b1010000000000100000010000001100001101000000000000000000000000000;
		8'd244: 64'b0100000000000110000000000000010000100000100000000000000000000000;
		8'd245: 64'b0010000000000000000000000000001000010000000000010001100000001000;
		8'd246: 64'b0000000000000100010000000000000000000000000000010000100000100000;
		8'd247: 64'b0000000000000000000100010000000000000000000000000000000000000001;
		8'd248: 64'b0000000001100100010000000000001000000000000000010000000000000001;
		8'd249: 64'b1110000011000110000000000010000000000000000000000000000000001000;
		8'd250: 64'b0100100000100000010001000000010000000000000000001000000000000000;
		8'd251: 64'b0101000000000000000000000101001000000000100100000010000000010100;
		8'd252: 64'b0010001000000000001000000000000000000000000000000001000000000000;
		8'd253: 64'b0000000000000001000000000000100000000000000000000000000010000000;
		8'd254: 64'b0000100001010000010000000010000010000000100000000001000001000000;
		8'd255: 64'b0000000000000001000100000000000000000000000000010000000101000100;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page1(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1000110010001011010000001000000000011100100100100001100001000000;
		8'd1: 64'b0010001010011000001010000000000000111000010100100000100011000000;
		8'd2: 64'b0000000000000000010000000111000001000000011100010010101000011101;
		8'd3: 64'b0001011010110010000001100001000000011001100011000010000100111001;
		8'd4: 64'b0101000000000001000011010000000011000000000000000000001011000000;
		8'd5: 64'b0000001000111000000010001100011000000000101100100000010000100001;
		8'd6: 64'b0001010011010100001001001100000000101000000000000000000001010001;
		8'd7: 64'b0000000111010100000001100001000000010000000010000100100111010000;
		8'd8: 64'b0101010000100011000000110010000100000100010100000001101000000010;
		8'd9: 64'b0100011000000000001000001000000100000000000000111000100010000000;
		8'd10: 64'b0111000100010000101001001101011010010100000010000000100000001000;
		8'd11: 64'b1001000001000001000000000010000000010001010100110010100000001011;
		8'd12: 64'b1010010001010001000000000000100000000011000100000010000000000010;
		8'd13: 64'b0000010000000010001000000000101000001011110010010011100000011010;
		8'd14: 64'b0100100000010010100010000100000011010000000000110000001000000101;
		8'd15: 64'b0110110000000001000101000000000110010000100000100010000010000000;
		8'd16: 64'b0010000011001100000000010001001011100000101111000100100000000001;
		8'd17: 64'b1010101000000000000000000101000100101000000001000011000001000000;
		8'd18: 64'b1000000110000000001111100000000000110000000000001000011000101000;
		8'd19: 64'b0100101000110011000010110100000010011010110100011000100000000000;
		8'd20: 64'b0010000000001001001000100000101100000001000001111000001001011010;
		8'd21: 64'b0011000111110000100010001011001110000111010000111000100010100101;
		8'd22: 64'b0000000001110010000001100000110001001000001010000000000001000001;
		8'd23: 64'b0011110000011000100000100000000000110101100010010010000100110000;
		8'd24: 64'b1000010100110010100100000011100000000101101001001000000110010011;
		8'd25: 64'b1010101010000001010000100101001110001111001100100010000000100000;
		8'd26: 64'b0001001010010101000001010000100001001011110000011000010000001001;
		8'd27: 64'b0000010110000100000000010000000000100000100000100100000100000010;
		8'd28: 64'b0100100000000010000100100000011100000001010010000000001010000010;
		8'd29: 64'b0110000010100001000100000000000010000000010000010111000010000000;
		8'd30: 64'b0100010010000001000000100000001000000000000001010000100000100000;
		8'd31: 64'b0000000100000010100000001110000000011000100001100100001011000000;
		8'd32: 64'b0100000001010000111000001001100000010000001100000000000000001000;
		8'd33: 64'b0001000000010101011001000010011000000000010100001110000000100000;
		8'd34: 64'b1001000100101000010000010100010100011000000101001000000001100111;
		8'd35: 64'b0000101110010010000001001000100100010000100000001000001010010001;
		8'd36: 64'b1100001001000000100101010100001100001001010000000100001000100001;
		8'd37: 64'b0110010110000001000101010000000000100011110000000001000010000101;
		8'd38: 64'b1000000001000101100100000001011000000100010011000010000000010100;
		8'd39: 64'b0000101010001000100010100001000000000010100010001100000000000000;
		8'd40: 64'b0110000100000100000001000011100010100000010001010000010001000000;
		8'd41: 64'b0000000101010100000000110010000000000100000010001001000000000010;
		8'd42: 64'b1000100100011000010000000000100000000010000000000110000100100000;
		8'd43: 64'b1001100110000100010010000100010010010000000001000101000101001100;
		8'd44: 64'b0101011000010101101101100001110001000110110100010001000000010000;
		8'd45: 64'b0000100010000001110000001001101100000010001100010100000010010010;
		8'd46: 64'b0000000000000000000000000000000100000100001000010100001111000000;
		8'd47: 64'b0100100100011101001010000000000000000000001001000010100010110000;
		8'd48: 64'b0011000000100000000100010001010001110000000000011000000001011001;
		8'd49: 64'b1000001100000001111010000000000000000010100100010000011000010100;
		8'd50: 64'b0000000010001111000000000100111100001101000101000011000100010000;
		8'd51: 64'b1010111010000011000011010000000000100100111000101010010000000000;
		8'd52: 64'b0111010000001000000100010010000000000010000001011000010000010000;
		8'd53: 64'b0100000000010100010000010000000000000000000000000011000000110000;
		8'd54: 64'b0100000000100000000000010101000000110001110001011010010001110001;
		8'd55: 64'b0000010001000110110000001100001000000000000000101100010000010000;
		8'd56: 64'b0000001100000001011001000000000001010000000010000101010011000001;
		8'd57: 64'b0100001000001000000001010110001100000010000011010100010001000100;
		8'd58: 64'b1000000001000011000000110000000000000010000101010010101000001101;
		8'd59: 64'b1000000000111000000110100000001000001000000010010011001101000011;
		8'd60: 64'b0001010100000000001001101010010111000011000000000010000010100100;
		8'd61: 64'b0000100000100001010100000101000011011110111000000101111100100100;
		8'd62: 64'b0010010010000110000001101000000001100010000001001111001000000000;
		8'd63: 64'b0000110000010000001001001011000000001100001000000001010000000000;
		8'd64: 64'b0100000101000001100010000001000100001100110000011000010000010011;
		8'd65: 64'b0000000101011000000010001101100110110000010100001000000010000000;
		8'd66: 64'b0001010000000010000000000000000000010000000000000011000100001000;
		8'd67: 64'b0000001100010000000101100001000001000100000100001010100010000110;
		8'd68: 64'b0000100001100010010000101011110001100000000100100100001001011000;
		8'd69: 64'b1000010000100100000000000010000000100110001101100010100000010010;
		8'd70: 64'b0000000000000000101101000010000000010000010101010100100000001000;
		8'd71: 64'b0011000110000100010110000000001010010011000000100001001100010100;
		8'd72: 64'b1010000100100111011000000001011010000000000100001000001000000010;
		8'd73: 64'b0000100000000000000001000100111000010100000000000000010011000000;
		8'd74: 64'b0111100000100000000000101000000100001110000000011101000001000001;
		8'd75: 64'b0001010010011100000000111100100001000000100001001000000000011000;
		8'd76: 64'b1000010000000010100101010001010100000101000110110001011000000000;
		8'd77: 64'b0100000100000000100010000100000100010000000101010000001110101000;
		8'd78: 64'b0010011010101110000001010100011100000000000010100110100000000010;
		8'd79: 64'b0101100000001110000010111000101001100000000011000000011000111001;
		8'd80: 64'b0100010000000101000001010010010001011000000100011000011101001100;
		8'd81: 64'b0001100010100000000000000000101010111100000001100000000010000001;
		8'd82: 64'b0100000000000000001000000000001000001100000000110111101000100000;
		8'd83: 64'b0000000100000101100101000100010101100011100000010001100100000000;
		8'd84: 64'b0000001010001000100000101110010010000000100000010001111001101000;
		8'd85: 64'b0000011000010001000000000000000000000100110001000000010000000000;
		8'd86: 64'b0010001101000000000011110000011010000010010101000000000101010101;
		8'd87: 64'b0001000011010010100000000001000000000001000110000000010000110101;
		8'd88: 64'b1000101010000010000010010000011100000000001000110000010100000000;
		8'd89: 64'b0001000000100100001000010010011010100010000000010100000100001010;
		8'd90: 64'b1100000001000110000010000000010011110000000010100001001000001001;
		8'd91: 64'b0001000000000010000110000010010000011001000000000001000010000001;
		8'd92: 64'b0000100100101010000000001001100000001011110010100010101010010010;
		8'd93: 64'b0000000110010011011010000001100000101000010100010000100011100010;
		8'd94: 64'b0010100000000001000010000011000001100000000001000000101100000000;
		8'd95: 64'b1000000100110001001100000000010000100000000000000100000000000000;
		8'd96: 64'b0000000110100000010110110010101000000000000001010010010011101100;
		8'd97: 64'b0001000100101000001100101011000000000001001010100010100000000001;
		8'd98: 64'b0010000000000010101000100001001101110010000000100100010000000010;
		8'd99: 64'b0000000110000110001000000100000110010000001000001010010000000000;
		8'd100: 64'b1001100100001001100100011000100101011101000000001001000010100100;
		8'd101: 64'b0011100100100000010000001110010101010000000001100100000100000100;
		8'd102: 64'b0100000000010100011110100000011001101000101001001000100000000010;
		8'd103: 64'b0001010001000000000010001010000000000011001000100100001000000010;
		8'd104: 64'b0000111000000000000100000000000000010010010000011111110001001001;
		8'd105: 64'b0010001000000011001100000000001000000000000000110010010000000000;
		8'd106: 64'b0000111000110000000010000001000000100100001100010000000011010001;
		8'd107: 64'b0000000010100001000001100001100010010001000000000000000000000000;
		8'd108: 64'b1000011100000000000100100000001000010001000011001100100100001000;
		8'd109: 64'b0100100010000100000010010010000001000000111000010000001100000111;
		8'd110: 64'b0010001000001010010000001010000001100100000111010101000001100000;
		8'd111: 64'b0011000010110100100010010000000001101010000010101000101000100000;
		8'd112: 64'b1101000001010000011100000001000000010000000001001110001000010000;
		8'd113: 64'b1001010000001000011000001000000010000010000001000001000100000000;
		8'd114: 64'b0101001000000010001100000010000000001100010101001101001001010010;
		8'd115: 64'b0010100000000101001001010010111100100001000000000010001010001111;
		8'd116: 64'b0000100000001001001101000001000111011000000000001001000100001001;
		8'd117: 64'b0000101100100011001000000010010100000100011001000000000001110011;
		8'd118: 64'b1010010100000000000001000110011000000100010000000010000000000100;
		8'd119: 64'b0000011001100100011000010000001110000011001011001100000000000010;
		8'd120: 64'b0011001010011001010101000000000011000000000100010000010000101010;
		8'd121: 64'b0000101001110100001110000000000101011000010100000000100100110000;
		8'd122: 64'b0000000100000000000110000000000010000001101110011001000000000010;
		8'd123: 64'b0000001000000000001000100000000000101010000000100000000000000000;
		8'd124: 64'b1100000001000100101001000001000011000100010001100000001010001011;
		8'd125: 64'b0001000010010010000000000000010010000000010000000000000000100000;
		8'd126: 64'b0000010000000011000100010001000000110110010001101000010000001000;
		8'd127: 64'b0100001000000110100000000010000000000010001100010000000000100010;
		8'd128: 64'b0100000000111000000111111001000001100110100010101100000101100101;
		8'd129: 64'b0001001110000010001000001100010100100000001001010010001101000000;
		8'd130: 64'b0000000101000101011010010000100000100001100001000101000100100000;
		8'd131: 64'b1000000000100000001001001000100010000000000001100100000100010000;
		8'd132: 64'b1110000010010010000010000110000010000000000000010000010000000110;
		8'd133: 64'b0100001010000001000100000001110000001001100001010001000000000110;
		8'd134: 64'b0011000000101001010001010001000000010010001001110000101001001100;
		8'd135: 64'b1100000000000000000000000100000000010000001001001011010011010000;
		8'd136: 64'b0000001100010000100010010000110010001010000001000000000010010101;
		8'd137: 64'b0000100100100010000000001001000001011000100110000000100100011000;
		8'd138: 64'b0011001100000100000000000100100000100001000011100000000100000100;
		8'd139: 64'b1000100000000100000001001000010010000101001000000010000101000100;
		8'd140: 64'b0011000010100100100100000100000000000000000000001100000000100000;
		8'd141: 64'b1001010010000001010000100110011011000000010000010000000010000000;
		8'd142: 64'b0000110010001000010010011010100000001000001100000000000000100000;
		8'd143: 64'b0010100000000000100000000011000110000010000000000000000000010100;
		8'd144: 64'b0000000010001001011000000010000010100101001010010001000000000100;
		8'd145: 64'b0100000000000000010011100010000100010001001010100000000000010000;
		8'd146: 64'b0000001000101000010001000000000010000000000000010010010001001000;
		8'd147: 64'b0100000000001000010000100011000011010010100000100000001110100101;
		8'd148: 64'b0000001001000010000000100000000001000001011010000000000000001000;
		8'd149: 64'b0000001101001100000100100100000010100000010010101000010001000001;
		8'd150: 64'b0010101000000110101000010010000010001011000010001010011000100010;
		8'd151: 64'b1010100000000101100001100000110100000000000000111100000000000001;
		8'd152: 64'b1010000000110001000000010000000000000000001000000001000001000000;
		8'd153: 64'b0000001000000000010000100010010010000010100100100001100101001010;
		8'd154: 64'b0000000010100010000101110100000110011011101010100001011000000000;
		8'd155: 64'b0001000110110100000000010010010010110001001101000001001100010000;
		8'd156: 64'b0000000010010010000010000000100000100000100100000000010000000110;
		8'd157: 64'b0010000100000010110010100000000000000000000000000010010010000100;
		8'd158: 64'b0011100000000010010000000000011010100000000101001000001000101010;
		8'd159: 64'b0011000110000110000100001000010010010010101100001000011000001000;
		8'd160: 64'b0000101001000100000010000011101000100000000000000010001000110010;
		8'd161: 64'b0000000000101000110100000010110000000110001001000000000000010000;
		8'd162: 64'b1001001010011000011100000100000001011000101001111000000010000010;
		8'd163: 64'b1000000100000101100000000000100100000001000000000010000100001000;
		8'd164: 64'b1100000100000110000000000000010010000100001011000000000110111100;
		8'd165: 64'b0000000000100110011100010000010100001000101001100000000100010000;
		8'd166: 64'b0000001100010110001100010100000010100001110100010011000001010010;
		8'd167: 64'b1100100000000000100101101001001011000100000000010010011001000010;
		8'd168: 64'b0111000010010001001000100110000000000000000001000000101101000000;
		8'd169: 64'b0010010110101000000000100000001000000001111000011100000000000000;
		8'd170: 64'b0100100000001001000000000011011111000011011110001001110010001010;
		8'd171: 64'b0010000000001011010000000010001100000100101000110001010001101011;
		8'd172: 64'b0001001000001000000000000000100000000000000000000000001000000000;
		8'd173: 64'b0001100000000100011000100000011000000000011000000000101010000100;
		8'd174: 64'b1001000110100010001110100000000100010001101000100001000010010000;
		8'd175: 64'b0101000010010000000000111000100001010000000000000101111010001000;
		8'd176: 64'b0100110001000100000110100001000000000010010110100010010000100101;
		8'd177: 64'b0100000000010101000000100100011010000000000010100011000001001001;
		8'd178: 64'b0100010000100000000101000000001000001000011010100000101100010011;
		8'd179: 64'b0000100101011010000100001010100100000000100010000000000000000010;
		8'd180: 64'b0010001011000000100101010000100000101010000001000100001000010000;
		8'd181: 64'b0010000101000001000000000001100000100000010000000110100010010000;
		8'd182: 64'b0100100100010001000001000000000000000011001110010010000000001101;
		8'd183: 64'b0010001111000000000000010100001000000010101010101000100101011000;
		8'd184: 64'b0000100011101001000010101011100001000000110001000001101000000000;
		8'd185: 64'b0000001101000001010101000001010000000100010100001001001100000000;
		8'd186: 64'b0001000100000010000011001100100000000100001000100010010000100000;
		8'd187: 64'b0000011110000000111100011000000000000001010000000000000000101010;
		8'd188: 64'b1001010010001010101000000001101000001000000000101010100100000101;
		8'd189: 64'b1010000000100000000000000000000000110000011001000000101011000100;
		8'd190: 64'b0000000100000001000000000001001000001001000011010000100010010000;
		8'd191: 64'b0001100001001000001001000111000000100011110011000000100101100110;
		8'd192: 64'b0100000000000001000001010110000011000110010000010001000001000000;
		8'd193: 64'b1100000001001011101010001000000011011101100000010000001000010110;
		8'd194: 64'b0100000010000100000101111000000001000011110001000010001000100001;
		8'd195: 64'b0100001110100000010000000100001011000011001000010100010000010000;
		8'd196: 64'b0100111000000000000101000001010100001000000001000010000100010110;
		8'd197: 64'b0010000001001101000000111001000001010000010000101001100100001010;
		8'd198: 64'b0000000001000000100001100001000101100000000010010001000000000000;
		8'd199: 64'b0000001011011011000010000110000010100100100100011100000010001100;
		8'd200: 64'b0001011000100100000001000000110110001000100101000000011100001000;
		8'd201: 64'b1000001110110000001000110000110000110000001001000011001000001011;
		8'd202: 64'b0000000000000100100000011000010100000000000000100000000010000000;
		8'd203: 64'b0000000010101100010100010000100000001000000111110001001001000000;
		8'd204: 64'b0000000110000000100001000010010010100001000000101010000000100010;
		8'd205: 64'b1001001010010000000000000000010011110000000100000000000100010100;
		8'd206: 64'b1000000000000000101011010000100100000000000000000000110001000010;
		8'd207: 64'b0110000000010011100100000111111010000000001100000101001101000011;
		8'd208: 64'b0100000000001000010000100000000001100000000000000100000001000000;
		8'd209: 64'b0110100000000100101000010010100000000000000010101010100110001000;
		8'd210: 64'b0001001100000001000110000010110101100010001001001000010000100000;
		8'd211: 64'b1011000000000000000001010110100000110000000000000010100001001100;
		8'd212: 64'b0000011110000000000000010110100001010100000000000100000001000000;
		8'd213: 64'b1001000000110000001000000110000010100011000000011001100001010100;
		8'd214: 64'b0001001111000000100000100001000000000110000000001000001100011000;
		8'd215: 64'b1010001001000000000010100000000100000000100000111000000110110000;
		8'd216: 64'b0001001000000000100001000000000000000010000000010001101000000100;
		8'd217: 64'b0111000001000000000100000010000000010000000000000011000001000001;
		8'd218: 64'b0010001000011000010000011010000000000000100100000000100111010001;
		8'd219: 64'b0010000000011000000000010000000000100001011100010100000000001000;
		8'd220: 64'b0001001000000010001100001000011100110001010000000000000110001100;
		8'd221: 64'b0000001010010000100100000000000010010011101000001000000101001001;
		8'd222: 64'b1000001000000000111110010010000100110100000100000000010000111111;
		8'd223: 64'b0000100010000100000000011100000000001001000100010100000011000000;
		8'd224: 64'b1000001000011100000010100010001011011000110000011000110001001010;
		8'd225: 64'b0000001000001000101000000000010010000100000000000101100000100100;
		8'd226: 64'b0110000001000000000010100100000001100001010000000001000011000100;
		8'd227: 64'b0000000011100000000100000010000000100101000000000000100000001001;
		8'd228: 64'b0000000000001000110000010101100011000100110001101000000000011100;
		8'd229: 64'b0000100000010000000010000001000000000000110100000001100100000000;
		8'd230: 64'b0000010100000100000000010000100000000101100000001110111001000000;
		8'd231: 64'b0000111100000000100001010000001010000010000100010000000010000000;
		8'd232: 64'b0000001010000010100001010000000000000000010100100000000001000100;
		8'd233: 64'b0110010100000010000000001000000000011101000010100101000001011100;
		8'd234: 64'b1001001000010011000000000010000000110100000000110100100100110001;
		8'd235: 64'b0100100100001000010100100000001001010000000100010000001010000000;
		8'd236: 64'b0000001001000000000100000010100000100100000001010000101100010000;
		8'd237: 64'b1010101011000000000000000000001100001000010001100100010000000000;
		8'd238: 64'b0100010000100000001000000001000000100111001010000110000000011000;
		8'd239: 64'b0100010010110010001100000000000100000001000100000000000000001101;
		8'd240: 64'b0000001000000000010100010101100100000000101000000000000001101001;
		8'd241: 64'b1000000001000100001001000001011000001000110001000000010000000100;
		8'd242: 64'b0010101010110000110001111000011100100010100010000000000000000001;
		8'd243: 64'b1011010000000101000010000001100011101000111000100000000000000000;
		8'd244: 64'b0100000100000110000000000100010100100010100000100000100010000000;
		8'd245: 64'b0010000000000100000010000001001010110100010000011011100010001000;
		8'd246: 64'b0100000100000100010000000000010000101000000000010000110010100000;
		8'd247: 64'b1100000000010001010100010000000100000001000000000000100000000001;
		8'd248: 64'b0000000001100101011110100000101000010000001010010000000000000001;
		8'd249: 64'b1110000111000110000000000010000010001000000000100100000000011000;
		8'd250: 64'b0100100100100000111001000000010010001000000000001000000000000000;
		8'd251: 64'b0101000010001100000000000101011000000000100100000010000000010100;
		8'd252: 64'b0011001000000010111000000000000000011000000100000011000000000101;
		8'd253: 64'b1000001000010001100000000100100000000000000001000000100010110000;
		8'd254: 64'b0100100001110000010000100010000010010000101000000001000001101000;
		8'd255: 64'b0000000010000001000100010001100001000000000000010100000101100100;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page2(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1101111011001011010000101100000000011110100100100001110001000000;
		8'd1: 64'b0010111010011100101010001000000011111000011100100000100011000000;
		8'd2: 64'b0000000000000010011001000111010001000000011110110010101000011101;
		8'd3: 64'b0011011011110011000101101001001000111001110111100010001110111001;
		8'd4: 64'b0101000000010001000111110010000011010000001000010000001111101000;
		8'd5: 64'b0000101010111000000010001100011000010000101100101000010011100001;
		8'd6: 64'b0001110011010101001001011100000110111100100001000001000101010001;
		8'd7: 64'b0010011111010100010011100001000000010001100110010101100111010000;
		8'd8: 64'b0101010000100011000000110110100101111100011100010001101000000010;
		8'd9: 64'b0100011000000110101000001000000101000000000001111000100010000100;
		8'd10: 64'b0111000100011000101101001101011010010100000011010011100000001100;
		8'd11: 64'b1001011001110001000010000011000000110001010100111111100100011111;
		8'd12: 64'b1010010001010101110000000100100000000111101100000111010001111010;
		8'd13: 64'b0000110011000010101000000001101000101111110010010011100110011010;
		8'd14: 64'b0101101000010110100010000100000011111100001000110010001000100101;
		8'd15: 64'b0110110000000001000101000000001111010110100001100110010011001001;
		8'd16: 64'b0010010011101110000000010011001011100100101111001101101000010001;
		8'd17: 64'b1110101100000010101001000101001100101000100001100011000001000000;
		8'd18: 64'b1010000110000000101111100000000000110010000010001000011000101000;
		8'd19: 64'b0101101010110111000111111100000010011010110100111001110010000000;
		8'd20: 64'b1010001000001001101000100101101100001001010001111001111111011010;
		8'd21: 64'b0011110111111000100011101011001111101111011100111010101010101101;
		8'd22: 64'b0000000001111010001001100110110001101000001010000000000001000001;
		8'd23: 64'b0011110010011000100000111010110010111101100010010010000110111000;
		8'd24: 64'b1000010110111110110100011011101000000101101001001000100110010111;
		8'd25: 64'b1010101010010101111010111111011110001111001100101110000101100101;
		8'd26: 64'b0001001010011101000001010000100101001011110001011000010010001111;
		8'd27: 64'b0010010110000101000000010000000000100001100000100100101101000010;
		8'd28: 64'b0100101100000010000100100000011110000011011110100000001110000110;
		8'd29: 64'b0110000011100001010100000010100010100001010011010111000110110000;
		8'd30: 64'b0100010010000001001100100000101110010000000001010000110001101000;
		8'd31: 64'b0001000100100010111000011110000101011000101001101100001011000000;
		8'd32: 64'b0100000101010000111000001001100010010000001110000000000000001000;
		8'd33: 64'b1001000001010101011001000110011000000100010101011110101100100000;
		8'd34: 64'b1001010100101010010000010110110100011010100101101100000001101111;
		8'd35: 64'b1010101111011010100001001000100110010000101011101000011110010001;
		8'd36: 64'b1101001101000010101101011111011110001011010010000100111001110101;
		8'd37: 64'b1110011110000001000111110001110001101011110000100001000010000101;
		8'd38: 64'b1000101001000101101101001101011001000100010011000010000000010110;
		8'd39: 64'b0011101110001100110011110001000100110011100010001101100000000001;
		8'd40: 64'b0110010100000110000011100111110011100000110001010100010011001100;
		8'd41: 64'b0011010101010100100110110011000000000100010010001001110000000010;
		8'd42: 64'b1000110101011010010001100001100000000010000100110110010100100010;
		8'd43: 64'b1001101110000101010010011111010010111000000001000101000101001100;
		8'd44: 64'b0101011000011101101101100001110001000111110100010001011101010110;
		8'd45: 64'b0010101110100001110011001001111100000011101100011100000010110011;
		8'd46: 64'b0000110100000100001000100000000100000100001000010100001111000000;
		8'd47: 64'b1110101100011101011011100100000000000000101001000110101011110100;
		8'd48: 64'b0011000000100001011100110001110011111000110010011110001111011001;
		8'd49: 64'b1100001110000011111010100001000001000010100100110000011100010101;
		8'd50: 64'b0000000110001111001000010100111100001101100101010011000100110010;
		8'd51: 64'b1010111010000011001011011000010010111101111000111010010001001110;
		8'd52: 64'b0111010001011010000101010010000110010110000001011100111110010000;
		8'd53: 64'b0101000100010100011101010000000000010000000010000011101001110000;
		8'd54: 64'b0100000111110111010000110101000001111011110111011010010001110001;
		8'd55: 64'b0010011011000111111000001111001000000100100000101100010010010000;
		8'd56: 64'b0100011100000001011111000001000001010000000111000101010011000001;
		8'd57: 64'b0110001000101100011001010110001101000010000111011100110001011100;
		8'd58: 64'b1000000001100011001000110000010001000011010101010110101001001101;
		8'd59: 64'b1000000000111000000110100101001001001100001010010011011101010011;
		8'd60: 64'b1001110110100101001001101010010111000111000000000010000110110101;
		8'd61: 64'b1000100100100001010101000111001011011111111001110101111100100101;
		8'd62: 64'b0110111011000110101001101000000001110010000001001111001101010000;
		8'd63: 64'b1000110010110100001001111011100001001100011000000011010011000000;
		8'd64: 64'b0100010101000011110010000001000100001101111100011100110000010011;
		8'd65: 64'b0110000101011000000110001111100110110000010101001000000010111001;
		8'd66: 64'b0101010000011010000000110001000000011000000010100011010101001110;
		8'd67: 64'b0000011100010101000111100101000001000110010101011010100010010110;
		8'd68: 64'b1000100001100010010001101111110011100111000101100100001001011000;
		8'd69: 64'b1000010000100110000100100010001000100110001101100010100100010010;
		8'd70: 64'b0000000001000000101101000010000110010100010101010100110000101000;
		8'd71: 64'b1011000110111100010110110001011010010111010011100101101100010100;
		8'd72: 64'b1010000100110111011000001001011010000000000100001100001010001010;
		8'd73: 64'b0000110011000100010011000100111100010100000000000001010011000000;
		8'd74: 64'b0111100001101000010000101000000100011110011000011101100101000011;
		8'd75: 64'b0001110010011100000001111110100001000000100111001000000010011000;
		8'd76: 64'b1000010001000010100101110001010100001101000111110001111000000001;
		8'd77: 64'b0100000100000010100010001100001100010100001111010010001111101000;
		8'd78: 64'b1010011011101110000001010101111100010000010010101110110000001011;
		8'd79: 64'b0101100000001111010010111010101001100000100011000000011000111011;
		8'd80: 64'b1110010100010101000001110111010001011000000100011100011101001101;
		8'd81: 64'b1101101010100100001000001000101010111100000001110010010110000001;
		8'd82: 64'b1100100100000000001100000000101000001100101000110111101100100010;
		8'd83: 64'b0010101100100101100101010110010101110011110001010001101101000000;
		8'd84: 64'b0011001010001000100000101110010110000010100001110011111001101000;
		8'd85: 64'b0001011100010001000001100101100000000101110001100011011100000000;
		8'd86: 64'b0011001101100000010011110000011010000010110101100000010101010101;
		8'd87: 64'b0001000011010011100100011001000000010001000110010001010000110101;
		8'd88: 64'b1000111011011010000010010100011110000110001010110000010101000000;
		8'd89: 64'b0011000000100101011000111010011110100011000000010100000100001010;
		8'd90: 64'b1101000001000110000010101000110111110000100111110011001100001111;
		8'd91: 64'b0001100000100110000110000010010100011001000000000001000010010011;
		8'd92: 64'b0000100110111010000010001101101000001011110010100010101010011010;
		8'd93: 64'b0100000110010011011010010001100101101000010100010000101011111010;
		8'd94: 64'b0010101000000101001010000111100001100010100001000000101101001000;
		8'd95: 64'b1100000101110001101100001000010001100000010001011111010000100100;
		8'd96: 64'b0010001110101001010110110010101100000000100001010010010111101100;
		8'd97: 64'b1001111100101000001110101011000010100001001010101111100000000101;
		8'd98: 64'b0010000000000010101000110001001101110011001100100100010000100010;
		8'd99: 64'b0111100111000110001000001101000110010000001001001110010011000000;
		8'd100: 64'b1001111100001001111100011000100111011101001000001101000110100100;
		8'd101: 64'b0011100100100000010000001110011101011000000001100100010100010100;
		8'd102: 64'b0101000011010110011110100101011101111000101001001100100000000110;
		8'd103: 64'b0101010101000011001010001010000010000011001000100110001000010010;
		8'd104: 64'b0000111100000001000100000000111110010010010010111111110001011011;
		8'd105: 64'b0010001000000111011101010000111000000000000000110010010000010010;
		8'd106: 64'b0000111100110000001010001001000000100111001100110000000011010001;
		8'd107: 64'b1001110010100001010001110001100010010001000010000000001001100000;
		8'd108: 64'b1001011100001000001100110010011000011001000011011110101100111000;
		8'd109: 64'b0100101010100100000010110010000011001010111000110100011100100111;
		8'd110: 64'b0110001000101011010000001010010001100100000111010101010001100100;
		8'd111: 64'b0011000010110100100010010001001011111010101011101000101101110000;
		8'd112: 64'b1101000001010011011100000011010000010000100101001110101000010000;
		8'd113: 64'b1001011000001000011111001000000010000010000011000011000110000000;
		8'd114: 64'b0101001000001010001100000010000000001101010101011111011001010011;
		8'd115: 64'b0010100000100101001101111110111100100001010001000010011111001111;
		8'd116: 64'b0000100110101001001101000001100111011001000001011011011100001001;
		8'd117: 64'b0111101100100011001010100010010101000100011001110000000001110011;
		8'd118: 64'b1010110100000010001011000111011001000110110010100010010000000100;
		8'd119: 64'b0000011101100100011000111000001110010111001011001101010000000010;
		8'd120: 64'b0011001011011111010101000000000111000010000110010000010001111010;
		8'd121: 64'b0100101111110111001110100000001111011100010110000000100100110001;
		8'd122: 64'b0000010110010101000110100000001010000011101110011001100101001011;
		8'd123: 64'b0011001001000000001100100000000000101010010000100000101100000000;
		8'd124: 64'b1100101001000100101001100001010011000100011001100010101011101011;
		8'd125: 64'b1011000010010010101000000100010010000000110000101001010010110000;
		8'd126: 64'b0110010001001011000101110001000000110110010001101001010000001010;
		8'd127: 64'b0110001010110110100000000010010100100010001101010100000000100110;
		8'd128: 64'b1100110000111010000111111111010001100110100010101100010111101101;
		8'd129: 64'b0001101111000111101000001110011111100000001001011110001101000010;
		8'd130: 64'b0100000111000111011011010000110100111001100001010101000111100111;
		8'd131: 64'b1000000000100010011001101000100010000000001011101100000100010000;
		8'd132: 64'b1110000010111011010010100110000010000100000000111000110001000110;
		8'd133: 64'b0100001010000001100110000001110100001011100101010101011111000110;
		8'd134: 64'b0011001000111011010001010101110100010010011001110000111001001100;
		8'd135: 64'b1100101000100100010100000100000100011000101001001111110111010000;
		8'd136: 64'b0001011100110000101110110000111011001011000111001010010110111111;
		8'd137: 64'b0000100100100111000000111001100001011001101110000000100100111000;
		8'd138: 64'b0011001100000100000000001100100000111001001011100010000100011100;
		8'd139: 64'b1001110000000110100011001000010110001101001001010010110101010100;
		8'd140: 64'b0011001010101100100100000100000100001000000000101100101011100011;
		8'd141: 64'b1001010010000001010000100110011011010110110000010000101010000100;
		8'd142: 64'b0100110010101000111110011010100000001000001111000000000000101000;
		8'd143: 64'b0010101000011000100000000011001110110011000000100000000000010111;
		8'd144: 64'b0000000010001001011001100110000010100101011110010001001000010100;
		8'd145: 64'b0100001000011000011011100011000100110001001010100110100001010000;
		8'd146: 64'b0000001000111101010001001000000111000000100010110011010001001111;
		8'd147: 64'b0110001001001000010010100011001111010010100011110100001110110101;
		8'd148: 64'b1100001101000010010000100000000001000001011010000000010000001001;
		8'd149: 64'b0010101101001110000100100110011110100111011011101000010001001111;
		8'd150: 64'b0010101010011110101100110110010010011011100010001010011000100010;
		8'd151: 64'b1010100000000101101001100000110110101010000010111100000100000001;
		8'd152: 64'b1110000000111011010001010011101000010101001101001001000001101010;
		8'd153: 64'b0000001000001000010100110010010010000011110110100001100101001010;
		8'd154: 64'b0001101110101010000101111111010110011111101111110001011010001000;
		8'd155: 64'b0001101110110110000001110011010011111011101101000001011100010101;
		8'd156: 64'b0000010010010010000110110000100000101000110100000000110000000110;
		8'd157: 64'b0010001100000010110010101000000010000000000000000010010010000100;
		8'd158: 64'b0011100000010010010001000100111010100010001101101000011000101011;
		8'd159: 64'b1111010110010110110100101000011110010110101101101000011000101000;
		8'd160: 64'b0011101101011110010010010111101001100000101000100110001011111011;
		8'd161: 64'b0001000000101000110100000010110010000110001011100001000000011000;
		8'd162: 64'b1011001110011001011101000100000001111000111001111110001010000011;
		8'd163: 64'b1000000100000101100110010000100101000001000000010010000100001000;
		8'd164: 64'b1101000100000110000100100000010010100100001011000000100110111100;
		8'd165: 64'b0000000000110110011101010010010100011000101011101001000100010010;
		8'd166: 64'b0000001100010110001100110111000010100101110111010011100101010111;
		8'd167: 64'b1101100001000000100101101001001111000100100000010110011001000010;
		8'd168: 64'b0111001010010001001000111110000000000001111001000100101101010011;
		8'd169: 64'b0010010110101010000110110000001000000001111001111100110000011010;
		8'd170: 64'b0110110000101101000000001011111111100111011110001001111010001010;
		8'd171: 64'b0010000000001011111000000010001101110100101000111001010011101011;
		8'd172: 64'b0001001000001010000000000110100100000100000000000001001000001000;
		8'd173: 64'b0001100100000100011010101011011000000010011000000000101010100110;
		8'd174: 64'b1001000110110110001110100000000100011001101001100101110011010001;
		8'd175: 64'b0101000010010000010000111000100001010000100000000101111010001000;
		8'd176: 64'b0100111101010100000110100011000100000010010110100110010000110101;
		8'd177: 64'b0100000001010101000001100100011110001000000010110011010001001001;
		8'd178: 64'b0100011000100000000111010110001001001000011010110000101101011011;
		8'd179: 64'b1000100101011010010110001010100100000000100110100000001000000110;
		8'd180: 64'b0010001011000000100101010000100000101010000101011111001101010100;
		8'd181: 64'b0010000101000001100000000001110000111000010001110110100010010000;
		8'd182: 64'b0100111101011001100001000001100100010011001110010010010000111101;
		8'd183: 64'b0010001111001000000000010100001001100010101010101110111101011000;
		8'd184: 64'b0100100011111001000110101011101001000001111001100011101110000000;
		8'd185: 64'b0001001101011001110101100001110000000110011101011001001100010001;
		8'd186: 64'b0001010101000010001011101100100000000100011000100010010100100100;
		8'd187: 64'b0001011110010000111110011001000100001001010110000000000100111010;
		8'd188: 64'b1011011010001010101010001001101000101010101001101011100110010111;
		8'd189: 64'b1110000101100000001000110100010001110001011001000100101111100100;
		8'd190: 64'b0100000100000001000100000001011100001001000011010100101010010010;
		8'd191: 64'b0001100101001000001001000111100101100011110011000100100101100110;
		8'd192: 64'b0100000001100001000011010110000111010110010000010001000001100000;
		8'd193: 64'b1100011001001011111010011001010011111111100000010000001101010111;
		8'd194: 64'b1110000010000100010101111001000001010011110001001011001000100001;
		8'd195: 64'b0101001110100010010001100111001011000011001100011101010000010010;
		8'd196: 64'b1110111010100100010101101011011100001110000001010010010101010110;
		8'd197: 64'b0111000001001101001010111001100101111000010110111001101100001110;
		8'd198: 64'b0000000001001101100011100001000101100010000010010011100000000000;
		8'd199: 64'b1010001011011011000010001110000010110100100100011100100010011100;
		8'd200: 64'b0001011000100100110101000010110111001000101111000100011100101001;
		8'd201: 64'b1000101110110010001000110010110100110010001101000011001000101011;
		8'd202: 64'b0000001000100100100000011100010111000000100000101010000110000000;
		8'd203: 64'b1000000110101101110110010010110000001000000111110001101001001010;
		8'd204: 64'b1000000110010110100001000010010010100011000000101010001000100010;
		8'd205: 64'b1001011011010000010001110000010011110110110100000100000100011101;
		8'd206: 64'b1100100000101000101011010100100100000010101001000000110001100110;
		8'd207: 64'b0110010101010011100100000111111010010000101100110111001101010011;
		8'd208: 64'b0101000000101000010000100011000001100000000010100100000001000100;
		8'd209: 64'b0110100000000111101000010010100001100000000010101010100110011000;
		8'd210: 64'b0001001100000011010110010010110101110010011001001001010100100000;
		8'd211: 64'b1011000000110000001001010110110100110000010010000010110101001100;
		8'd212: 64'b0000011111000000000110010110100001010101001000010100000001000110;
		8'd213: 64'b1011000000110001011000000110010010110011000000011001101001010100;
		8'd214: 64'b1001111111000000100100110001110100010110010000001010101100111100;
		8'd215: 64'b1110001111000000000010110000001110000001100000111000000110110001;
		8'd216: 64'b0111001000000101110001100000000100000010000010111001101001000110;
		8'd217: 64'b0111000001000000000100000010000000010011010000000011010001000001;
		8'd218: 64'b0010001011011000011000011010011010000001110100000010100111010001;
		8'd219: 64'b0010000000011000100100010011000100100101011100010100011100011000;
		8'd220: 64'b0101001000001110101101011000011101110011010101000010000110001100;
		8'd221: 64'b0000001111111000101100110001000010010011101110001000000101001001;
		8'd222: 64'b1000011000100000111111010010010100111100100100000000110000111111;
		8'd223: 64'b0000101110000111001001111100000011001001100100010100000011100000;
		8'd224: 64'b1000011010011100000010101110001011011100110000011000110001101010;
		8'd225: 64'b1010101000101001101000000000110010100100001010011101100000101100;
		8'd226: 64'b0110000101000100010110101100000101100001010000000001000111100100;
		8'd227: 64'b0010011011100000000101010010110101111101001000000010101100001001;
		8'd228: 64'b0000000000001000110000110101100011000100110011101000101100011100;
		8'd229: 64'b0100100000011000010010010101001000110001110101000001100100000100;
		8'd230: 64'b0100111111000100101000110001100000000101110000011110111001010001;
		8'd231: 64'b1000111100010000110001010100001010000011010100011000010010000000;
		8'd232: 64'b0000001010000010100101010010010000000010010100100000010001010101;
		8'd233: 64'b1110011101000010000000001000001001011111001010100111000001011100;
		8'd234: 64'b1011011010010011000010001010000000110100100100111110100100110011;
		8'd235: 64'b0110100100111000010110100001001101110100000100010011001010000100;
		8'd236: 64'b0000001001000001100100101010100000100100000001010100101100011000;
		8'd237: 64'b1010111011010111001011011000001100001011110001101101011000010100;
		8'd238: 64'b1100011011100000001000000001100101100111001111000110110000011000;
		8'd239: 64'b0101011010110011101100000000100110100001001100000000000000111111;
		8'd240: 64'b0110101000000010010100010101100100000010111010000000000111101001;
		8'd241: 64'b1110001001000100101001000001011010001000110011011010010000011100;
		8'd242: 64'b0010101010110000110001111100011110100010110010001000010011001001;
		8'd243: 64'b1011010000010101000010000001100011101000111001110001010010010000;
		8'd244: 64'b0100101101000110000000001100010100100011100001100000101010011010;
		8'd245: 64'b0010000010100100000010010011001010110100110000011011100010001000;
		8'd246: 64'b0100110100001100010000000000010000101100001000110000110010111010;
		8'd247: 64'b1100100100010001010110110010000100000001010010000010100000110001;
		8'd248: 64'b1100000001100101011110100000101001010001101010010010100001001001;
		8'd249: 64'b1110000111010110000001000010000011001000000000100100011000011011;
		8'd250: 64'b0111100100101110111001100001111110001001000010001001010000000100;
		8'd251: 64'b0101000010001100000101100101011000001100110111110111110000010110;
		8'd252: 64'b1011001000000010111000001000010101011010000100000011100010000101;
		8'd253: 64'b1000001000010001100010010100110000010001001001000001100011110100;
		8'd254: 64'b0111101111110000011010100011000010010000111110010001000101111000;
		8'd255: 64'b0000000010000001000100010001100001000001000100010101010101100101;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page3(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1111111011011011111101101100000010111110100110111001111011001000;
		8'd1: 64'b0010111010111110101010011010001011111010111100100010100111000010;
		8'd2: 64'b0010010000000010111011100111010001100010011110110110101100011111;
		8'd3: 64'b1011011011110011000101101001001000111001110111100010001110111001;
		8'd4: 64'b1101000001010011000111111110100011010001101000010100101111101000;
		8'd5: 64'b0000101010111000000110011100011000111000101110101000010011100111;
		8'd6: 64'b0101110011010101101001111110000110111100100001010101010101010001;
		8'd7: 64'b1011011111010100011011100001000000110001100110010101101111010001;
		8'd8: 64'b0101011100100011000010110110100101111100111100010101101000000010;
		8'd9: 64'b0101011010000110101110001000001101000010100011111100100010000100;
		8'd10: 64'b1111000110011000101111001101011010110100000011010011100001001100;
		8'd11: 64'b1001111001110001000111000011000000110001011101111111100110011111;
		8'd12: 64'b1010010001010111110001100101100001000111101100001111010101111010;
		8'd13: 64'b0010110011000010101000001001101000101111110010010011100110011010;
		8'd14: 64'b0101101010010110101010000111001011111100011100110110001010100101;
		8'd15: 64'b0110110100000011011101001010001111010111100001101110010011001011;
		8'd16: 64'b0010010011101110000000011111001111100100101111001101101000010001;
		8'd17: 64'b1110101101100011101001000101001110101000100001100011000001000100;
		8'd18: 64'b1010000110001000111111100100000000111010000010001100011000101000;
		8'd19: 64'b0101101010110111101111111100001011011010110100111001110110100001;
		8'd20: 64'b1010101000011101101011101101101101101011010101111011111111011010;
		8'd21: 64'b0011110111111011110011101011001111101111111110111010111110111101;
		8'd22: 64'b0000100001111010001001100110110001101000011110000000000001101001;
		8'd23: 64'b1011110010011000100000111011110110111101101010010010000110111001;
		8'd24: 64'b1000010110111111110100011011111100000101101001101000100111010111;
		8'd25: 64'b1110101010010101111010111111011110001111011101101110000101110101;
		8'd26: 64'b0001001010011101000001011100110101001111110101111000010010011111;
		8'd27: 64'b0010010110011101010000010010000100100101100000100100111111000110;
		8'd28: 64'b0100101100100010100110100000011110100011011110100000001110000110;
		8'd29: 64'b0110011111100001011100000010110010100001010111011111000111110010;
		8'd30: 64'b0100010010000001001100100100101110010000000001010001110001101001;
		8'd31: 64'b0001001100100110111110111110001101111100101001101100011111001100;
		8'd32: 64'b0100000101011000111000001101100010010000011110000001000010011000;
		8'd33: 64'b1001000101010101011001000110011100000100011101011110101100101110;
		8'd34: 64'b1001010110111010110000110110110100011010101101101110000001101111;
		8'd35: 64'b1011101111111011101001101001110110010000101111111001011110010001;
		8'd36: 64'b1101001101010011101101011111111110011011010010110100111001111111;
		8'd37: 64'b1110011111000011010111111101111011101011110000101001001010010101;
		8'd38: 64'b1100101001001101101111001111111001001101010011001010000011010110;
		8'd39: 64'b1011101111001100111111110001000100110011100010001101101100000001;
		8'd40: 64'b0110010100010110000011101111110011100000110111010100010011001100;
		8'd41: 64'b0011010101010100100111110011001000000100010110001001110000000010;
		8'd42: 64'b1000110101011011010001100001101010000010010100110110010100100110;
		8'd43: 64'b1001101110000101110110011111010010111000000101000101000101011100;
		8'd44: 64'b1111011100011101101101111011110001010111110100110011011111010110;
		8'd45: 64'b0010101111110011110011011001111111000011101110011100011111110011;
		8'd46: 64'b0000110100000100001100111101010100000101001000010100001111000100;
		8'd47: 64'b1110101100011101011011100100000011000000101001100110111011110100;
		8'd48: 64'b0011101110100001011111111001110011111000110010111110111111111101;
		8'd49: 64'b1110101110000011111011100011010011000010100100110000011100010111;
		8'd50: 64'b1000100110001111001000110100111100001101101101010011000100110011;
		8'd51: 64'b1010111010100111001011011001011010111101111000111011010001001111;
		8'd52: 64'b0111010001011110100101010010001110010110000001011100111110010011;
		8'd53: 64'b0101000100010100011101010000000000010000100110000011101001110000;
		8'd54: 64'b0101000111110111010100110101100001111011110111011010010001110001;
		8'd55: 64'b0010011011000111111001001111001010000100100001101100010110110010;
		8'd56: 64'b0100011101000101011111000001000111010101100111000101110011011001;
		8'd57: 64'b0110001100111111011101110110011101100010010111111100111001011100;
		8'd58: 64'b1110000001100011001001110000010001000011010101010110111011001101;
		8'd59: 64'b1000010000111000100111110101001011001100101010010011011111010111;
		8'd60: 64'b1001110110100101001001101010010111001111100001000010011110110101;
		8'd61: 64'b1100100100110001110101000111111011011111111101110101111101100101;
		8'd62: 64'b0110111011000110101001101000000001111010000001101111001101010101;
		8'd63: 64'b1000110010110100011101111011110001101100111110000011011011100110;
		8'd64: 64'b0100010111000011110010000001000100001101111111011101110001110011;
		8'd65: 64'b0111100111011000100110001111100110110010010101011000101010111001;
		8'd66: 64'b0101111010011010010000110111001000011000101010100011010111011111;
		8'd67: 64'b1110011100010111000111100101010101100110010101111110110110010110;
		8'd68: 64'b1001100001100010010101101111110011110111000101101100011011011110;
		8'd69: 64'b1100010100111110000100110010001011100111001101100010101100010010;
		8'd70: 64'b0001010111000100101111000111000110011100110101010100110000101000;
		8'd71: 64'b1011111110111101011110110001011011010111010111100101101110111100;
		8'd72: 64'b1010000100110111011000101001011010000001000100001100001010001110;
		8'd73: 64'b0000110111000101111011000100111100011100010000001011010011000100;
		8'd74: 64'b1111100101101001110001111000000110111110111100011111110101011111;
		8'd75: 64'b0001110010011100000111111110100001000000100111001000100010011111;
		8'd76: 64'b1000110001000010100111110011010101111101100111110001111111011001;
		8'd77: 64'b0110010100001010100010001100111100010100001111010010111111101100;
		8'd78: 64'b1010011011101111000001010101111100010001010010101111110100001011;
		8'd79: 64'b0111100000001111110011111011101001100000101011000000011000111011;
		8'd80: 64'b1111010100110101010011110111010101011100010111011100011111101101;
		8'd81: 64'b1101111010100100101000001100101010111100000001111011010110000001;
		8'd82: 64'b1100100101000000001100000000101011001100111000110111101100101010;
		8'd83: 64'b1010101101100111100111010110010101110011110001110001101111000100;
		8'd84: 64'b1011001010001100100001111110011110110110100001111011111011101100;
		8'd85: 64'b0101011100010001100111110111101100000101110001100011011110010000;
		8'd86: 64'b1011001101100000010011110001011111010010111101101100010101110101;
		8'd87: 64'b1001000011010011100110111001000010010001010110010001010110110101;
		8'd88: 64'b1000111011011110000111010101011110000110101011110000110101000001;
		8'd89: 64'b0011101100100101111000111010011110100111001100110100000100011010;
		8'd90: 64'b1111000001000110000010101100110111110100101111110011011100001111;
		8'd91: 64'b0001100000101110000110000011010100011001001000000001000010010111;
		8'd92: 64'b0000100110111010011011001101101000001111110010101010101011011010;
		8'd93: 64'b0100110110011011011010011001100101101001110100110010101111111010;
		8'd94: 64'b0110101110001101001010010111100001111110100001000100111101001000;
		8'd95: 64'b1101010101110001111100101000110011100000110101011111111000100100;
		8'd96: 64'b0010001110101001010110110010101100001001111111010011010111101100;
		8'd97: 64'b1001111110101010111110101011100010100111001010101111110000000101;
		8'd98: 64'b1110001000010011101001110001001101110011001100100110010000100010;
		8'd99: 64'b0111110111100110011000101101000110010001001101001110010011100000;
		8'd100: 64'b1001111100001001111100011000100111011101001100001101000110100100;
		8'd101: 64'b0011100100100000010001001110011101011000001001100100010110010100;
		8'd102: 64'b0101000011011110011110111101011101111100101111001100111001010111;
		8'd103: 64'b0111011101000011001010001010000010010011011000100110001110010010;
		8'd104: 64'b0000111110001001101100010000111111010010010010111111110001111011;
		8'd105: 64'b0010001000000111011101110000111100000101000101110010010100111010;
		8'd106: 64'b0000111110110011001111001001100110101111001100110000011111010001;
		8'd107: 64'b1011110110110001010001110011100010010001000010000010001001100000;
		8'd108: 64'b1111111100101110001100110010011000011111000011011110111100111000;
		8'd109: 64'b0101101010100110000110111011000011001010111001110100011100100111;
		8'd110: 64'b0110011001101111010000001010010101100100001111010111010011100100;
		8'd111: 64'b0111000110110101101010010011001111111011101011101000101101110000;
		8'd112: 64'b1101000001010011011101100011010010010000110101001110101001110100;
		8'd113: 64'b1001011000001110011111001100100010010010000011000011111110000000;
		8'd114: 64'b0101001000001011001100010010000110011101010111011111011001010011;
		8'd115: 64'b0110100000100101001111111110111101100101110001000010111111101111;
		8'd116: 64'b1000110110101011101111010001100111011001000001011011011100101001;
		8'd117: 64'b0111101100101011001010101010010101001100011001110010100011110011;
		8'd118: 64'b1010110111000010001011001111011001000110110011100010010000000100;
		8'd119: 64'b0101011101110100111000111000001111010111011111001101010000000010;
		8'd120: 64'b0011001111011111010101000000000111000010010110110000010001111010;
		8'd121: 64'b0101101111110111001110100000001111011110010111000000100100111001;
		8'd122: 64'b1000010110010101100110100001001010010011111110011001100101001011;
		8'd123: 64'b0011001001010010001100100000000000101010010100100100101101000000;
		8'd124: 64'b1100101001000100101001110001010011001100011011100010101011101011;
		8'd125: 64'b1011000010010011101000001100010010000000110011101001010010110010;
		8'd126: 64'b0111010001001011000101110001101000110110010001101001011000001010;
		8'd127: 64'b0111001010110110100000011010010100100110101101010100000000100111;
		8'd128: 64'b1100110000111010010111111111010001100110110010101100110111101101;
		8'd129: 64'b0111101111000111111011001110011111101010001011111110011101000110;
		8'd130: 64'b1100000111000111011011111000110100111001100001010101110111100111;
		8'd131: 64'b1000000010110010011001101001100011000010101011111100010110010010;
		8'd132: 64'b1110000110111011010010100110001110000101010000111000110001000110;
		8'd133: 64'b0100001010000011100111000101110101001011110101010111111111000111;
		8'd134: 64'b1011001010111011111001010101110100110010011011110001111111011101;
		8'd135: 64'b1100111000110100111100010101000110111000101001001111110111010010;
		8'd136: 64'b0011011100110000101110110001111011001011000111111010110110111111;
		8'd137: 64'b1001100100110111000010111101100101011001101110101100110100111001;
		8'd138: 64'b0011001100100110000000001100110000111001001011100010100100111100;
		8'd139: 64'b1001111000001110100011001000010110001101001011011010110101010100;
		8'd140: 64'b0111101010101100100101000100100100001010010000101100111011100011;
		8'd141: 64'b1001010010000001010100101110011011010110110001010000111010001100;
		8'd142: 64'b1100110010101000111110011010101010011001001111000000000000101010;
		8'd143: 64'b0010101000111010101000000011001110110011010000100010001001010111;
		8'd144: 64'b0000000110001001011001110110100110100111011110010101101100111100;
		8'd145: 64'b0100001000111001011111110011001100110001001010100110100001110010;
		8'd146: 64'b0000101000111111111001001000100111000000100010111011010001001111;
		8'd147: 64'b0111001001001100010010101011101111010010111011110100011110110111;
		8'd148: 64'b1100001101000010010000100000000001011001011010000000010001001101;
		8'd149: 64'b0010111101001111000111100110011110100111111011101000010011001111;
		8'd150: 64'b1010111010011110101101110110011010011011100010001010111000101010;
		8'd151: 64'b1010101000011101101011101000110110101010000011111100000100001001;
		8'd152: 64'b1110000100111011011011011011101000011101001111001101101001101010;
		8'd153: 64'b1000001000001000010100111010011011010011111111100111110101001010;
		8'd154: 64'b0001101110101010100101111111111110011111101111111001111110101000;
		8'd155: 64'b1001101110110111001101111011010011111011101101010001011100010101;
		8'd156: 64'b1000011010010110000110110010110000101010110110000000110100001110;
		8'd157: 64'b0010001110000010110011101000010010010000000001001010110010000100;
		8'd158: 64'b0011110000010011011001100100111110100010001101101010011000101011;
		8'd159: 64'b1111011110110110110100101001011110010110101101101010011000101010;
		8'd160: 64'b0011101101111110010010010111101001110001111000100111001011111011;
		8'd161: 64'b0001100100101000110101000010110010010110001011100001001000011100;
		8'd162: 64'b1011101110111111011101011100001001111100111001111110101010000111;
		8'd163: 64'b1001000100100101100110010000101101000001100000010010100101001001;
		8'd164: 64'b1111100100100111101100110000010010111100001011000000100110111100;
		8'd165: 64'b0000000000110110011101110010010100011000101011101001000100010011;
		8'd166: 64'b0010001101010111001100110111000010100101110111010011110101010111;
		8'd167: 64'b1101100001000000110101101011011111000110110000010110011011000010;
		8'd168: 64'b0111001010110001001000111111000000100101111001000100101101010011;
		8'd169: 64'b1010010110101010000110111010001000000001111001111100110001011010;
		8'd170: 64'b0110110010101111100000001011111111101111111111101001111010001010;
		8'd171: 64'b0010001000101011111000001010101101110101101000111001011111101011;
		8'd172: 64'b0001011000001010000000001110101100100100010110000001001100001000;
		8'd173: 64'b0011100100000100011010111011011000010011011001110010101011100110;
		8'd174: 64'b1101100110111110001110100001000101011001101001100101111011010011;
		8'd175: 64'b0101000010010000010001111000100001011000100000100101111010101010;
		8'd176: 64'b0100111101010110010110100011000101000010010110100110010010110101;
		8'd177: 64'b0100100001010111101001100100011110001100010010111011110001001001;
		8'd178: 64'b0100011001100010000111110110001001001001011010110001101101111011;
		8'd179: 64'b1011100101011010010110001010110100100000110110100100001000000111;
		8'd180: 64'b0010011011000000101101011000100100101010000101011111101101010101;
		8'd181: 64'b0010000101000101110000010101110000111001010001110110100010010000;
		8'd182: 64'b0100111101011001100001000011100100011011011110010010010100111101;
		8'd183: 64'b0011001111101000011000110100101111100011101010101110111101011010;
		8'd184: 64'b0100100111111101000110101011101011001001111001100011101110000010;
		8'd185: 64'b1001001101011001110101101101110100010110011111111011001100010101;
		8'd186: 64'b0001010101000010001111101101100000000100011000101111010101100100;
		8'd187: 64'b0001011110011000111110011001000110011101010110000011000100111011;
		8'd188: 64'b1011111010001010101010001001101010101110101001101011100110010111;
		8'd189: 64'b1110000101100000001110110110010001110001011001000100101111100100;
		8'd190: 64'b0100001101000011000100000001011100001011000011010100101010010010;
		8'd191: 64'b0001100101101100011001000111101101110011110011000110100101110110;
		8'd192: 64'b0100011101100101000011010110000111110110010000110001000111100000;
		8'd193: 64'b1100011001001011111010011011010011111111100010010110001101110111;
		8'd194: 64'b1110101010000100011101111001110101010011110001001011011011110001;
		8'd195: 64'b1101011110100111010001110111011011000011111100011101011010010110;
		8'd196: 64'b1110111010101100010101101011011100111110001001010010010101110110;
		8'd197: 64'b1111000001001101001010111011100111111000010110111001101100011110;
		8'd198: 64'b0000010001001101101011101001000101110010000011010011100000000000;
		8'd199: 64'b1010001011011011000010001110100010111101100111111100100011011100;
		8'd200: 64'b0001011000110100110101000010110111001000101111011100011100101001;
		8'd201: 64'b1010101110111110001100110010110100111010001101000011001000101011;
		8'd202: 64'b0000001110100101110100011101110111001010100001111011000110000100;
		8'd203: 64'b1000101110101111110110010010111100101000100111110001101111001010;
		8'd204: 64'b1000000110110110100001001111110010101011011000101010011000100110;
		8'd205: 64'b1011011011011000011101110001011011110110110101110100000110011101;
		8'd206: 64'b1110100000101010101011011101110100101010111011001000110001101110;
		8'd207: 64'b0110010101010011111110000111111010010001111100110111101101110111;
		8'd208: 64'b0101000000101000010010100011011001101100010110100100000001000110;
		8'd209: 64'b0110100000101111111000010010100001100000100010101010100110111000;
		8'd210: 64'b0001011101000011010111010010110101110111011001101001110101100000;
		8'd211: 64'b1011010000111100001001010111110110110000010110000110111101001100;
		8'd212: 64'b0000011111100000000110011110100011010101011000010100000001000110;
		8'd213: 64'b1011000100110001011111100110010010110011001101011011101001010100;
		8'd214: 64'b1001111111100010100110110101111110010110010011101110101100111110;
		8'd215: 64'b1110001111001100000010110000001111000001100100111000000110110001;
		8'd216: 64'b0111011000000111110001110000010100000110000010111011101001100110;
		8'd217: 64'b1111001001001010011100000010001001010011010000000111010011000001;
		8'd218: 64'b0010001111011001111100011011011010000001110100001110110111010101;
		8'd219: 64'b1010001100111001100100010011100100100101011100011100011100011100;
		8'd220: 64'b0111001001001110101101011110011101110011010101000111000110001110;
		8'd221: 64'b0000001111111001101100110001000011010011111110001101000101001001;
		8'd222: 64'b1000011000100001111111010010010100111100100100010000110110111111;
		8'd223: 64'b0000101110000111001011111100000011001001100100010100001011100000;
		8'd224: 64'b1100111010011100100011101110001011111110111001011010111001101010;
		8'd225: 64'b1010101010101011101000000000110010101100001010011111100010101110;
		8'd226: 64'b0110000101000100010110101100000101111101010000101001001111100110;
		8'd227: 64'b0010011111100000011101110010110101111101001010000010101100101011;
		8'd228: 64'b0100010010001001110001110101111011100100110111101000111100111100;
		8'd229: 64'b0101101100011000010010010101001000110001110111000001100110010110;
		8'd230: 64'b0101111111011100101001110101100000011101110110011110111001010001;
		8'd231: 64'b1000111100011001110001010100001010010011010100011001010010000000;
		8'd232: 64'b0001001110001010110101010110110000000010010110101100010011010111;
		8'd233: 64'b1111111101001010010001111000011001011111001010100111000001111100;
		8'd234: 64'b1111011010010011100010001110000100110100111100111110100100110011;
		8'd235: 64'b0111110100111000011110100001001101110100010100010111011011000100;
		8'd236: 64'b0010001101000011100110101011100000100110000001010100101100111000;
		8'd237: 64'b1010111111010111101011011000001110001011110101101101011000010111;
		8'd238: 64'b1100011011110000001000000101110111100111001111001110110011111000;
		8'd239: 64'b0101011010110011101100001010110110100001001100000000000000111111;
		8'd240: 64'b1110101110100011010101010111110101000010111010000000000111101101;
		8'd241: 64'b1110101101000111111001000001011011111000110011011010010000011100;
		8'd242: 64'b0010101010111000110001111100011110100010110010101010010011001101;
		8'd243: 64'b1111011010010101001010101001100111101000111101110001010010110000;
		8'd244: 64'b0100101101000110000000101111110100100011100001110000101010111010;
		8'd245: 64'b0010000010100101000010011111011010110101111001011011100010001000;
		8'd246: 64'b0100110100001100010000001001110000111100011000110100110111111111;
		8'd247: 64'b1100100100010001010110110010000100000001011110010010100001110101;
		8'd248: 64'b1111010001101101011110100010101001010101101110011011100011001101;
		8'd249: 64'b1110000111010110010001000010000011001010010000100101011010111011;
		8'd250: 64'b0111100100111110111011100001111111011101100010001001010000000101;
		8'd251: 64'b0101100010001111000101100101011010001100110111110111110000010110;
		8'd252: 64'b1011001000110010111010001000010111011010000100100011100010000111;
		8'd253: 64'b1000011000011101110010010101110111010001001001001001100011111110;
		8'd254: 64'b0111101111111001011010101111011010010100111110010011001101111000;
		8'd255: 64'b0000000010000101000101010111100001000001001110010101010101100101;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page4(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1111111111011011111101101101001010111110100110111011111011001000;
		8'd1: 64'b0010111010111110101010011010001011111010111100100010100111000110;
		8'd2: 64'b0011011000000010111011100111010001100011011111110110101100111111;
		8'd3: 64'b1011011011110011000101101001101000111001110111111011001110111001;
		8'd4: 64'b1101000101110011000111111110100011010001111000010111111111101000;
		8'd5: 64'b0101101011111010110110011101011000111000101110101000111011100111;
		8'd6: 64'b0101110011010101101001111110000110111100100011010101010111010001;
		8'd7: 64'b1011011111010100011011100001000000111001100110011101101111010101;
		8'd8: 64'b0101011100100011000010110110100101111111111100010101111100001010;
		8'd9: 64'b0101011110000110101110101000001101000010100011111100100010011100;
		8'd10: 64'b1111100110011000101111001111111010110101001011010011100001001100;
		8'd11: 64'b1001111001110001000111010011010000110001011101111111100110011111;
		8'd12: 64'b1010010001110111110001100101101001000111101101001111011101111010;
		8'd13: 64'b1110110011100110101100011101101000101111110010010011100110011010;
		8'd14: 64'b0101101011010110101010100111001011111110011101110110001011100101;
		8'd15: 64'b0110110100100011011101001010001111110111100101101110010011001011;
		8'd16: 64'b1010010011101111101000111111001111100101101111011101101100010001;
		8'd17: 64'b1110101111100011101001000101001111111000100001100011010001000100;
		8'd18: 64'b1010001110001000111111100110000000111010000010001110011000101000;
		8'd19: 64'b0101111010111111101111111101101011011110110100111011110110100011;
		8'd20: 64'b1010101000011101101011101111101101101011111101111011111111011110;
		8'd21: 64'b0011110111111011111011101011101111101111111110111010111111111111;
		8'd22: 64'b0100100011111010011001100110110001101001011110000011000001101001;
		8'd23: 64'b1011111010011000100001111011110110111101111010010010100110111011;
		8'd24: 64'b1010010110111111110100011011111110001101101101101010100111010111;
		8'd25: 64'b1111111110110101111110111111011110101111011101111110000101110101;
		8'd26: 64'b0001001010011111000001111110110111001111110101111000010010011111;
		8'd27: 64'b0010010111011101010010010010000100100101110010110100111111000111;
		8'd28: 64'b1100101100110010101110100001011110100011111110100000001110000110;
		8'd29: 64'b0110011111101001111101010010111110100001010111011111000111111110;
		8'd30: 64'b0101010010000001001101100100101110010000010001010001110001101001;
		8'd31: 64'b0001101110100110111110111110011101111110101001101101111111101100;
		8'd32: 64'b0100000101111000111000001101100011010001111111100001110111011000;
		8'd33: 64'b1011000101010111011001000110011100100100011101011110101100101110;
		8'd34: 64'b1001010110111010110100110110111100111010101111101110000001101111;
		8'd35: 64'b1011101111111011101011101001110110111000101111111011011110010001;
		8'd36: 64'b1101001101010011101101011111111110011011011010110110111101111111;
		8'd37: 64'b1110011111000011110111111101111011101011110000101011001010010101;
		8'd38: 64'b1100101011001111111111001111111001001101010011001111000011010110;
		8'd39: 64'b1011101111001100111111110001100100110011100010011101101100000001;
		8'd40: 64'b1110110101111110011011101111110011101100110111010100010011111100;
		8'd41: 64'b0011010101010110100111110011001010010100010111001001110000000010;
		8'd42: 64'b1100111101011011011001100001101010000011010100111110010101100111;
		8'd43: 64'b1001101110000101110110011111010010111000101101000101000101011100;
		8'd44: 64'b1111011110011101111101111011110001010111110100110011011111010110;
		8'd45: 64'b0110101111110011110011011001111111000011101110011100011111110011;
		8'd46: 64'b0000110100000100011100111101010100001101001001010100101111100100;
		8'd47: 64'b1110101100011101011011100100100011001000101001100110111011110100;
		8'd48: 64'b1011111110100101011111111001110111111010110010111110111111111101;
		8'd49: 64'b1110101110010011111011100011010011000010100100110100011100110111;
		8'd50: 64'b1000100110001111001000111100111101001101101101011011010101110111;
		8'd51: 64'b1111111010100111101011111001011010111101111000111111110011001111;
		8'd52: 64'b0111010011011110100101010010001110010111000001111100111110010011;
		8'd53: 64'b0101000100010100111101110001110000110000110110000011101011110001;
		8'd54: 64'b1101000111110111110100110101110001111011111111011011011001111001;
		8'd55: 64'b0110011011000111111001001111001010010110111001101100010111110010;
		8'd56: 64'b0100111101000101011111010101000111010101100111000111110011111001;
		8'd57: 64'b0110001101111111011101110110011101100011010111111100111001011100;
		8'd58: 64'b1110001001100011011101110100010011010011010101110110111011001101;
		8'd59: 64'b1010010000111001101111110101001111001110101010010011011111010111;
		8'd60: 64'b1001111110100101001011111010010111001111100001011010011111111101;
		8'd61: 64'b1100110100110101110101000111111011011111111101110111111101100111;
		8'd62: 64'b0110111011000110101001101000000001111010000001101111001101010111;
		8'd63: 64'b1000110010110100011101111011110001111100111110000011111011101110;
		8'd64: 64'b0100010111101111110010000001010100001101111111011101110001111011;
		8'd65: 64'b0111100111011001100110001111100110110011010101011000101010111001;
		8'd66: 64'b0101111110111010010100110111001000111010101010100111010111111111;
		8'd67: 64'b1111111100010111000111110101010101100110010101111111110110010110;
		8'd68: 64'b1001100001100010010111101111110111110111000101101100011011011111;
		8'd69: 64'b1100011101111110000101110111001011100111101101100010101100010010;
		8'd70: 64'b0001110111000100101111000111000110111101110101010100110000101010;
		8'd71: 64'b1011111110111101011110110001011011110111010111100101101110111100;
		8'd72: 64'b1110000100110111011000111001011010000101000100001100001110001110;
		8'd73: 64'b0000110111000101111011000100111100011101010011011011010011000100;
		8'd74: 64'b1111110101111001110001111000001111111111111100011111110101011111;
		8'd75: 64'b0001110011011100010111111110100001000000100111001000100011011111;
		8'd76: 64'b1100110101010110100111111011110111111101110111110001111111111001;
		8'd77: 64'b0110010100011011100010001100111100010100001111010010111111101101;
		8'd78: 64'b1010011111101111100111110111111100010101010010101111110101001011;
		8'd79: 64'b0111100010001111110011111011101001100101101011000000011000111011;
		8'd80: 64'b1111010101110101010111110111110101011100011111011101011111101101;
		8'd81: 64'b1101111010100110101000001100101010111100100011111011010110001001;
		8'd82: 64'b1100100101000000001100000000101011001100111000110111101100101010;
		8'd83: 64'b1010101101100111100111010110010101111011110001110001101111000100;
		8'd84: 64'b1011001010001100100001111110011110110110110001111011111011101100;
		8'd85: 64'b0101011100010001100111110111101100000101110001110011011110010001;
		8'd86: 64'b1011001101100100010011110111011111110110111101101100011101110101;
		8'd87: 64'b1001000011110011100110111001000010010001110110010001011110110101;
		8'd88: 64'b1000111011011111100111010101011110001110101111110000110111001001;
		8'd89: 64'b1011101100100101111000111011111110110111001100111110000101011010;
		8'd90: 64'b1111000011000111111010101100110111111100111111110011011100101111;
		8'd91: 64'b0011100000101110000110000011010100011001001000000001000010010111;
		8'd92: 64'b0000101110111010011011001111101000001111110111101010101011111011;
		8'd93: 64'b0100110110011011011010011111110111101101110110110010101111111010;
		8'd94: 64'b0110101111001101011010010111100001111110100011000100111101101000;
		8'd95: 64'b1101010101110001111100101000110011110000110101011111111000101100;
		8'd96: 64'b0010011110101001111110111110111100101001111111010011111111101100;
		8'd97: 64'b1001111110101010111110101011100010100111001010101111111000000101;
		8'd98: 64'b1110001000010011101001111001101101110011001100100111010000100111;
		8'd99: 64'b0111110111110111011001101101000111010101001101001110010011100100;
		8'd100: 64'b1101111100001001111101011010101111011101001100001101000110111100;
		8'd101: 64'b0011100100100000010001001110011101011001101001100101010110010110;
		8'd102: 64'b0101100011011110011111111111011111111110101111011101111001010111;
		8'd103: 64'b0111011101000011001010111010000011010011011110100110001111010010;
		8'd104: 64'b0110111110001001101100011000111111010011011010111111110111111011;
		8'd105: 64'b0010001001000111011101110000111100001101000101110011110100111011;
		8'd106: 64'b0010111110110011011111101001101110101111011100110010111111011001;
		8'd107: 64'b1011110110110001010001110011100010010001001010000010001001100001;
		8'd108: 64'b1111111100101110011101110110011001011111000011111110111101111111;
		8'd109: 64'b0101101010100110000111111011000011001010111001110100011100100111;
		8'd110: 64'b0110011001101111010001001010110101101100001111010111010011100101;
		8'd111: 64'b0111000110111101101010010111011111111011101011101000101101110000;
		8'd112: 64'b1101000001010011011111100011010010110000110101101111101001110100;
		8'd113: 64'b1001011000001110111111001100100110010011000011000011111110100000;
		8'd114: 64'b1101001000011011001100010010000110011101010111011111011001011011;
		8'd115: 64'b0111100001100101001111111110111101100101111001000010111111101111;
		8'd116: 64'b1000110110101011101111010001100111011101000001011011111100111001;
		8'd117: 64'b0111101100101011101010111010011101001100011001110010100011110011;
		8'd118: 64'b1110110111010010001011001111011001010110110011100010010001000100;
		8'd119: 64'b0101011101110100111100111000001111010111011111001101010001000010;
		8'd120: 64'b0111001111111111010101000110000111100011010111110000010001111111;
		8'd121: 64'b0101101111111111001110100001001111011110011111000001100100111001;
		8'd122: 64'b1011010110010101100110101001101010010011111110111001100101011011;
		8'd123: 64'b0011001001010010001100100000000001101010010100100100101111000010;
		8'd124: 64'b1100101001000100111001111001010011001100011011111010101011101011;
		8'd125: 64'b1011000010111011101000001100110010100000110111101001010010111010;
		8'd126: 64'b0111011001001011001111110001101010110110010001101001011000011010;
		8'd127: 64'b0111101010110111100010111010110100100110101101010101000100100111;
		8'd128: 64'b1100110000111011110111111111010001100110111010111100110111111101;
		8'd129: 64'b0111101111000111111011001110011111101010001011111110011101000110;
		8'd130: 64'b1100000111000111011011111000110110111101100001010101110111100111;
		8'd131: 64'b1000001010110010011001101001100011000110101011111110010110010010;
		8'd132: 64'b1111000110111011010011100110001110000101011011111000111001000110;
		8'd133: 64'b0100001010000011110111001111110101001011110111010111111111011111;
		8'd134: 64'b1011011011111111111001010101110100110010011011110101111111011111;
		8'd135: 64'b1100111000110100111100010101000110111000101001001111110111010010;
		8'd136: 64'b0011011110111001101110111011111111101111000111111010110110111111;
		8'd137: 64'b1001100100111111010010111111100101011001101110101100110100111001;
		8'd138: 64'b0011101100110110001000001100110000111001101011100010100100111100;
		8'd139: 64'b1001111000001110100011001000010110001101001011011010110101010101;
		8'd140: 64'b0111101011101100100101000101101100001010010000101101111011100011;
		8'd141: 64'b1001010010000001010100101110111011010110110001010000111010001100;
		8'd142: 64'b1101111010101000111110111010101010011101101111000010100010101010;
		8'd143: 64'b0110101000111010101000000011001111110011010010100010001001010111;
		8'd144: 64'b0100000110001001011001110110100110100111011110010101101100111100;
		8'd145: 64'b0100101000111001011111110011001100110011001010101111100001110010;
		8'd146: 64'b1010101110111111111101001100101111000001100110111011010001001111;
		8'd147: 64'b0111001001001101010010101111101111010111111111110100011110110111;
		8'd148: 64'b1100001101000010010000100001000001011001011010000000010101011101;
		8'd149: 64'b0010111101101111010111100110011110100111111011101001011011001111;
		8'd150: 64'b1010111010011110101111110110011010111011100010001010111010111110;
		8'd151: 64'b1010101010011111101011101000110110101010000011111100000110001011;
		8'd152: 64'b1111010100111011011011111011101000011101001111001111101001111010;
		8'd153: 64'b1000001010001000010100111010011011110011111111100111110101101010;
		8'd154: 64'b0001101110101010100111111111111110011111101111111001111110101001;
		8'd155: 64'b1101101110110111011101111011010111111011101101010011011110010101;
		8'd156: 64'b1000011010011110100110110010110000101010110110000000110110001110;
		8'd157: 64'b0010101110001010110011101010011110010000001001101110110110000100;
		8'd158: 64'b0011110000010111011001100101111110100010001101101010011000101011;
		8'd159: 64'b1111011110110110110100101001011110010110111101111010011010101010;
		8'd160: 64'b0011101101111110010010010111101101110001111001100111001011111011;
		8'd161: 64'b0101100110101000110101000010110010010111001011110001001000011100;
		8'd162: 64'b1011101110111111011101011100001101111110111101111110101010100111;
		8'd163: 64'b1001000100100101100110010000101111100001101000011010100101001101;
		8'd164: 64'b1111100100100111101100111010010010111110101011000000100110111100;
		8'd165: 64'b0000000000110110011101110010110100011000101011101001000100011111;
		8'd166: 64'b0010001101010111001100110111001110100101111111010011110101010111;
		8'd167: 64'b1101100111000000110101101111011111010110110000011111011011000011;
		8'd168: 64'b0111001011110101001000111111000000100101111001000110111101010011;
		8'd169: 64'b1010010110111010000110111010001000000001111001111100110101111010;
		8'd170: 64'b0110110011101111100000001111111111101111111111101001111010001010;
		8'd171: 64'b0010001110111011111001001010101101110101101010111101011111101011;
		8'd172: 64'b0101011100001010000100001110101101100100010110011001111100101000;
		8'd173: 64'b0011110100000101011010111011011000110011111001110010101011110110;
		8'd174: 64'b1101100111111110001111100101111111111001101101101101111011010011;
		8'd175: 64'b0101001010010000010001111100100001011000101100100101111110101010;
		8'd176: 64'b0100111101010110010110100011011101000010010110100111111010110101;
		8'd177: 64'b0100100001010111101001100100011110001100010010111011110001101001;
		8'd178: 64'b0100011101100011000111110110001011001011011010110101111101111011;
		8'd179: 64'b1011111111011110010110001010110110100000110110100100001000000111;
		8'd180: 64'b0010011011000010101101111001101100101010000101011111111101010101;
		8'd181: 64'b0010000101000101110000010101110110111101011001110110100011010000;
		8'd182: 64'b0100111101111001100001010011101100011011011110010010110110111101;
		8'd183: 64'b0011001111101010011100110100101111101011101010101111111101111010;
		8'd184: 64'b1100101111111101000110111011101011001101111001101011101110000010;
		8'd185: 64'b1001001101111001110101101111110100110111011111111011101110010101;
		8'd186: 64'b0001010101000010011111101111100000000100111001101111010111110100;
		8'd187: 64'b0001011110011000111110011001000110011111010111010011100100111011;
		8'd188: 64'b1011111010101010101010001101101010111111101001101011100110110111;
		8'd189: 64'b1110101101100010001110110110011101110001011001000101101111100100;
		8'd190: 64'b0100001101010011000100000001011101001011000011010100101110010010;
		8'd191: 64'b0101100101101100011001000111111101110011111011000111100101110110;
		8'd192: 64'b0100011101100101000011010110100111111111010000110001100111100000;
		8'd193: 64'b1110011001001011111010011011010011111111100010110111001101110111;
		8'd194: 64'b1110101010000100011101111001110101011111110001001111111011111011;
		8'd195: 64'b1101011110100111010001111111011111000011111100011101011010010110;
		8'd196: 64'b1110111010101100011101101011011100111110001001110010110111110111;
		8'd197: 64'b1111000001001101001010111011110111111000010111111001101100011110;
		8'd198: 64'b0011010001001101101011101011000101110010000011110011100010100000;
		8'd199: 64'b1010001011011011000011001110110110111101100111111100100011011110;
		8'd200: 64'b0001111101110100110101010010110111001000101111011100011100101001;
		8'd201: 64'b1010101110111110001100110010110100111011001111000011001000101011;
		8'd202: 64'b0000001110100101110101011101111111001110100001111011000110000101;
		8'd203: 64'b1010101110101111110110111010111110101000101111110001101111001010;
		8'd204: 64'b1000000110110110101001001111110010101011111101101010011000100110;
		8'd205: 64'b1111011011011000111101110001011011110110110101110100000110011101;
		8'd206: 64'b1110100010101010101011011101110100111011111011001010111011101110;
		8'd207: 64'b0110010101010011111110010111111110010001111100110111101101110111;
		8'd208: 64'b0101001000101010010010100011011011101100010110101101101001000110;
		8'd209: 64'b0110100010101111111000010010100001100000100010101010100110111000;
		8'd210: 64'b0001011111000011010111110110111111110111011001101001110101100000;
		8'd211: 64'b1111010010111100101101010111110110110000010110100110111101001100;
		8'd212: 64'b0000011111100000001111011110100011110111011000010100001001000110;
		8'd213: 64'b1011000100110011011111100111010010110011001101011011101001110100;
		8'd214: 64'b1001111111101010100110110101111110110110011011101110101101111110;
		8'd215: 64'b1110001111001100000010111000001111001101110101111000000110110001;
		8'd216: 64'b0111011000000111111001110000010100000110000010111011111101100110;
		8'd217: 64'b1111001001001010011100000010001001010011010000000111010011000001;
		8'd218: 64'b0010001111011001111110011011011010110001110101001111110111010101;
		8'd219: 64'b1010101101111001100100010011101100100101011100011100011100011101;
		8'd220: 64'b0111011011001110101101011110011101110111010101000111000110001110;
		8'd221: 64'b0000101111111001101100111001000011011011111110001101000101011001;
		8'd222: 64'b1000011000100001111111010010010100111100100100010000110110111111;
		8'd223: 64'b1111101110010111001011111100000011001001110101110100111011100001;
		8'd224: 64'b1100111010111100101011101110001011111110111101011110111001111010;
		8'd225: 64'b1010101010101011101000000010110010101101001010111111100010111110;
		8'd226: 64'b0111000101000100010110111100010101111101010100101001001111100110;
		8'd227: 64'b0010011111101000011101110010110101111101001010000011101100101011;
		8'd228: 64'b1100010010001001110001110101111011100100110111101000111100111100;
		8'd229: 64'b0101101101011000010110010101001001110001110111000001100110010110;
		8'd230: 64'b1101111111011100101011110101101000011101110110011111111011110001;
		8'd231: 64'b1000111110011001110101010100001010011011010100011001111110000001;
		8'd232: 64'b0001011110011010110101010111110100000010010110101101010011010111;
		8'd233: 64'b1111111101001010010001111010011001011111001010100111000001111110;
		8'd234: 64'b1111011010011011100010001110001110110100111100111110100100110011;
		8'd235: 64'b0111110100111000011110100001001101110100010100011111011011000100;
		8'd236: 64'b0010101101000011100110101011101010100110000011011101101100111000;
		8'd237: 64'b1010111111010111101011011000001110001011110101101101011000010111;
		8'd238: 64'b1100111011110000001100000101110111100111001111001111110011111000;
		8'd239: 64'b0111011010110011101100001110111111100001001100000000010000111111;
		8'd240: 64'b1111101111100111111101010111110101000010111011001100000111111101;
		8'd241: 64'b1110111101000111111001000101011011111000110011111110010000011100;
		8'd242: 64'b0011101010111000110001111100011110100010110010111010010011001101;
		8'd243: 64'b1111011011010101001010101011100111101000111101110001010010110001;
		8'd244: 64'b0110101101001110000000101111110100100011100001110010101010111110;
		8'd245: 64'b0010000010100101001010011111011010111101111001011011100011001000;
		8'd246: 64'b0100110100001100010010001101110001111100011000110100110111111111;
		8'd247: 64'b1100100100110101010110110010001100000011011110010010100001110101;
		8'd248: 64'b1111110001101101011110110011101001010101101110011011100011001101;
		8'd249: 64'b1110000111010110110001100010000011001010010000100101011110111011;
		8'd250: 64'b0111101100111110111011100001111111111101100010001101110100101101;
		8'd251: 64'b0101100010001111000101100101011010001110110111110111111001010110;
		8'd252: 64'b1011001000110010111110001000010111011010000100100011100110000111;
		8'd253: 64'b1000011000011101110010010101110111110001011101001001100011111110;
		8'd254: 64'b0111101111111001011010101111011010010100111110010011001101111000;
		8'd255: 64'b0001000010010101000101010111100011000001011110010101010101110101;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page5(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1111111111011011111101111101001110111110110110111011111011001000;
		8'd1: 64'b0110111010111110101010011010001011111010111100100010100111100110;
		8'd2: 64'b0011011000100010111011100111111001101011011111110110101100111111;
		8'd3: 64'b1011011011110011001101101001101010111001110111111011001111111101;
		8'd4: 64'b1101001101110011000111111110100111010001111010010111111111101000;
		8'd5: 64'b0101101011111110110110011101011110111010101110101001111111100111;
		8'd6: 64'b0101110111011101101101111110100110111100110011010111010111010101;
		8'd7: 64'b1011111111010101011011111001000111111011100110011101101111010101;
		8'd8: 64'b0101011100111011100110110110101101111111111100010101111100111011;
		8'd9: 64'b0101011110000110101110101000011111000010100011111100101010011100;
		8'd10: 64'b1111110110011000111111001111111110110111001011010011100101101100;
		8'd11: 64'b1001111101110001000111010011011000110101011101111111100110011111;
		8'd12: 64'b1010110101110111111001100111101001100111101101001111011101111010;
		8'd13: 64'b1110111011100110111100011101101000111111110010011011100110111010;
		8'd14: 64'b1101101011010110101010100111011111111110011101111110101011110101;
		8'd15: 64'b0110111100100011111101001010001111110111101101111110010111001011;
		8'd16: 64'b1010011011111111101001111111001111110111111111011101101111010001;
		8'd17: 64'b1110101111100111101001000101011111111010100001100011011001000111;
		8'd18: 64'b1010011110001001111111100110001000111011001010001110011000101000;
		8'd19: 64'b0101111010111111101111111111101111011110111110111011110110101011;
		8'd20: 64'b1010111110011101101111101111101101101111111101111011111111011111;
		8'd21: 64'b1011111111111011111111111111101111101111111110111011111111111111;
		8'd22: 64'b0100100111111010011101100110110001101101011110000011000001101001;
		8'd23: 64'b1011111010011010100011111011110111111111111010011110101110111011;
		8'd24: 64'b1011010111111111110110011011111110001101101101101111100111010111;
		8'd25: 64'b1111111111110111111110111111011110101111111101111110000101110101;
		8'd26: 64'b0001001010011111000001111111111111001111110111111000010010011111;
		8'd27: 64'b0010010111011111011010010010000100100101110011110101111111000111;
		8'd28: 64'b1100101100110010101110100001111110101011111111101000001111100110;
		8'd29: 64'b0111011111101001111101011111111111100001011111011111000111111110;
		8'd30: 64'b0101110010000011001101100100101111110000010001010001110001111001;
		8'd31: 64'b0001101110101110111110111110011101111110101001101101111111111100;
		8'd32: 64'b0101001101111100111100011101100011010011111111111001110111011000;
		8'd33: 64'b1011001101110111011001001110011100100101011101011110101101101110;
		8'd34: 64'b1011010110111110110100110110111100111010101111101111000001111111;
		8'd35: 64'b1011101111111011101111101001110110111100101111111011111110010001;
		8'd36: 64'b1101001101110011111111111111111110011111011110110110111101111111;
		8'd37: 64'b1110111111000011110111111111111011111011110010111111001111010111;
		8'd38: 64'b1100101011101111111111001111111011101111110011101111100111011110;
		8'd39: 64'b1011101111101100111111110001100100110011100010011111111100100001;
		8'd40: 64'b1110110101111110011011101111110011101100110111010100110011111100;
		8'd41: 64'b0011010101011110100111110011001010010100010111001001110000000010;
		8'd42: 64'b1100111101011011111001100101111011000111010100111110010101100111;
		8'd43: 64'b1101101110110101110110011111010110111000101101001101010101011100;
		8'd44: 64'b1111011111011101111101111011111011010111110101110011011111111110;
		8'd45: 64'b1110101111110011110011011001111111000111101110011100111111110111;
		8'd46: 64'b0000110100000100011101111111110100001101001001010100101111101100;
		8'd47: 64'b1110101101011101111011101100110011001100101101100110111011110100;
		8'd48: 64'b1111111111101111011111111101110111111010111011111110111111111111;
		8'd49: 64'b1110101110010011111011100011010111100010110100110110011100110111;
		8'd50: 64'b1000100110001111001000111100111101101101101111011011010101111111;
		8'd51: 64'b1111111010100111101011111001011010111101111011111111110011001111;
		8'd52: 64'b1111010011011110100101010111001111010111000001111100111110010111;
		8'd53: 64'b0101000100010100111101111001110000110000110110000011111011110101;
		8'd54: 64'b1111001111110111111100110101110101111011111111011111011001111001;
		8'd55: 64'b1110011011000111111001001111011010010110111101101100011111110011;
		8'd56: 64'b0100111101010101011111010111000111110101100111000111110111111011;
		8'd57: 64'b0110101101111111011101110110011101100011010111111110111001011100;
		8'd58: 64'b1110001011101111011101110100010011110111011101110110111011001101;
		8'd59: 64'b1010010000111001101111110101011111011110101110011011011111011111;
		8'd60: 64'b1101111110100101011011111011010111001111100001011010011111111101;
		8'd61: 64'b1101110100111101110111010111111111011111111101111111111111110111;
		8'd62: 64'b0111111011000110101101101001001011111010010001101111001101110111;
		8'd63: 64'b1010110011110100011101111011110001111110111110001111111111101110;
		8'd64: 64'b0100010111111111110111000001010100001101111111011101110001111011;
		8'd65: 64'b1111100111111101100110001111100110110111110101111010101010111001;
		8'd66: 64'b0101111110111010011100110111111000111010101010100111010111111111;
		8'd67: 64'b1111111100010111001111110111010101101110011101111111110110010111;
		8'd68: 64'b1011101001100110011111101111110111111111000111101100011111011111;
		8'd69: 64'b1100011101111110110101110111001011101111101101100010101100010010;
		8'd70: 64'b1001111111100100111111000111000110111101110101010101110000101011;
		8'd71: 64'b1011111110111101011110110001011011110111010111100101101110111100;
		8'd72: 64'b1110000100110111111000111001111010000101000100011100011110001110;
		8'd73: 64'b0000110111001101111011001100111110011101110011011111110011000100;
		8'd74: 64'b1111110101111001110011111100101111111111111100011111110101011111;
		8'd75: 64'b0001110011111100010111111111100001000000100111001001100011011111;
		8'd76: 64'b1100110101011110100111111011111111111101110111110001111111111001;
		8'd77: 64'b0110010100011011100010001100111100011100011111010011111111111101;
		8'd78: 64'b1010011111111111100111110111111100010101010010101111110101011011;
		8'd79: 64'b0111100010001111110011111011101101100101101011010101011010111111;
		8'd80: 64'b1111010101110101010111110111110101011100011111011101011111101101;
		8'd81: 64'b1111111010100110101011111101101011111100100011111011010110001001;
		8'd82: 64'b1100100101100000001100000000101011011101111000110111101100101010;
		8'd83: 64'b1110101101100111100111010110010101111011110001110001101111000100;
		8'd84: 64'b1011001010001100100101111110011110110110110001111011111011101111;
		8'd85: 64'b1101011100010101100111110111101100000111110001110011011111010011;
		8'd86: 64'b1011101101110110110011110111011111110111111111101111011101110101;
		8'd87: 64'b1001000011110011110110111001000110011001110110011011011110111101;
		8'd88: 64'b1000111111011111100111011101011110001110101111111000110111001001;
		8'd89: 64'b1111101110110101111100111011111110110111001100111110000101011010;
		8'd90: 64'b1111000111000111111110101101110111111100111111110111011101101111;
		8'd91: 64'b0111100000101110000111000011010100011001011001000001000010110111;
		8'd92: 64'b1110101111111010011011101111101100001111110111101010101111111011;
		8'd93: 64'b0100111110011011011110011111110111101101110111110010101111111111;
		8'd94: 64'b0110101111001101011110011111101001111111111011000100111101101000;
		8'd95: 64'b1101010101110101111100101000111111110001110101011111111001101100;
		8'd96: 64'b0010011111101001111110111110111100111101111111110011111111101101;
		8'd97: 64'b1001111110101010111110101011100010100111101010101111111001100101;
		8'd98: 64'b1110001000010011101011111001101101110011001100100111011000110111;
		8'd99: 64'b0111110111110111011001101101000111010101001101001110010111100100;
		8'd100: 64'b1101111100011001111111011110101111011101001110001101000110111100;
		8'd101: 64'b0011100100100000010001001111011101011011101001110101011110010110;
		8'd102: 64'b0101110011011111111111111111111111111110111111111101111001010111;
		8'd103: 64'b0111011101000011001010111010001011110011011110100110001111010110;
		8'd104: 64'b1110111110001011101100011000111111010011011010111111110111111011;
		8'd105: 64'b0010011011000111011101110010111100101111001101110111110100111011;
		8'd106: 64'b1010111110111011011111101011111110101111011100110010111111011001;
		8'd107: 64'b1011110110111001010011110111100010010011001110010010011001100001;
		8'd108: 64'b1111111100101111011101110110011011011111010011111111111101111111;
		8'd109: 64'b0101101010100110000111111111011011001010111001110110011100110111;
		8'd110: 64'b0110011001111111010001011010110101101101001111010111011011100101;
		8'd111: 64'b0111001110111101111010010111011111111011101011101100111101110110;
		8'd112: 64'b1101100001010111111111100011010010110100110101111111111011110101;
		8'd113: 64'b1001011000001110111111001110100110110011000011001011111110101000;
		8'd114: 64'b1101001000011011001100110010000110011101010111011111011001111011;
		8'd115: 64'b0111100111100101011111111110111101110111111001000010111111111111;
		8'd116: 64'b1011111110101011101111010011100111011101000001011011111100111001;
		8'd117: 64'b0111101100101011101010111110111101001100111001111010111011110111;
		8'd118: 64'b1110111111010111001011001111011001010111110011100010111001000100;
		8'd119: 64'b0111011101111101111100111000001111010111011111001101010101000011;
		8'd120: 64'b0111001111111111110101010111001111100111011111110000011001111111;
		8'd121: 64'b0101101111111111001110100001001111011110011111000001100100111101;
		8'd122: 64'b1011010110011101100110101001101010010011111110111001101101011011;
		8'd123: 64'b0011001001010010001100100000000101101111010101100110101111001010;
		8'd124: 64'b1100101001001100111001111001010011001100011011111010101011101011;
		8'd125: 64'b1011010010111011101010001100110010100100110111101001010110111011;
		8'd126: 64'b0111011001001011001111110001101010110111010001111011011010011010;
		8'd127: 64'b0111111110110111100010111010110100100110111101010101000101100111;
		8'd128: 64'b1100110001111111110111111111010011101111111011111110111111111111;
		8'd129: 64'b1111101111001111111011101110111111111010111011111110011101011110;
		8'd130: 64'b1101000111000111011011111000110111111101100011110101111111100111;
		8'd131: 64'b1100001010110010011001101101100011010111111011111110111110010010;
		8'd132: 64'b1111000110111011110011100110011111000111011111111000111001100110;
		8'd133: 64'b0100001010000111111111001111110101001011110111110111111111011111;
		8'd134: 64'b1011011011111111111101010101110101110011011011110101111111011111;
		8'd135: 64'b1100111010110100111100111101100110111010101011001111110111010010;
		8'd136: 64'b0011111110111101101111111011111111101111000111111011110111111111;
		8'd137: 64'b1001100100111111010010111111110101011001101110101100110100111011;
		8'd138: 64'b0011101100110110001010001101110000111001101011100010100100111100;
		8'd139: 64'b1001111000001110100111101000010110011101011011011110111101111101;
		8'd140: 64'b0111101011101110100101000101101100101010010100101101111011110111;
		8'd141: 64'b1001010011000001010100111110111011110110110001010000111010001100;
		8'd142: 64'b1101111010101110111111111010101010011111101111000011100010101010;
		8'd143: 64'b0111101000111010101101000011001111110011010010100010001001010111;
		8'd144: 64'b0100100110001001011001110110100110100111011110010101101100111110;
		8'd145: 64'b0101101000111011111111111011001100110011001110101111100101110011;
		8'd146: 64'b1011101111111111111101001101101111000001100110111011011001001111;
		8'd147: 64'b0111011101101111010110101111111111110111111111110100111110111111;
		8'd148: 64'b1100001101101010010000111011000001011001011010000000010101011111;
		8'd149: 64'b1110111101101111010111100110011111100111111011101101011011001111;
		8'd150: 64'b1010111010011110101111111110111010111011111010001010111011111110;
		8'd151: 64'b1010111010011111101011101000110110101010100011111110100110001011;
		8'd152: 64'b1111010101111011011011111011101000111101001111111111101101111010;
		8'd153: 64'b1011001011001000010100111010011011110011111111100111111101101010;
		8'd154: 64'b0101111111101110100111111111111110011111101111111001111110111101;
		8'd155: 64'b1101101110110111111101111011110111111011101101010011011110110101;
		8'd156: 64'b1010111010011110100110111110110100101010110110000000110111001110;
		8'd157: 64'b0010101110001011110011101010011110010000001001111110110110000100;
		8'd158: 64'b0111111000011111011001110111111110100010001101101010011000101111;
		8'd159: 64'b1111011110110111110101101001011110110110111101111010011010101011;
		8'd160: 64'b0111101101111110111010111111111101111101111101101111001011111011;
		8'd161: 64'b0111100110111000111101100010110011011111101011111001001100011100;
		8'd162: 64'b1111101111111111011101011100011101111111111101111110101010100111;
		8'd163: 64'b1001000101110101101110011000101111101001101010011110100101001101;
		8'd164: 64'b1111101110101111101100111010110010111111101011000010100111111100;
		8'd165: 64'b0000010000110110011101110010111100011000101011101001001110011111;
		8'd166: 64'b1011001101010111001100110111001110100101111111110011110101010111;
		8'd167: 64'b1101101111100011111101101111011111010111110000011111011011000111;
		8'd168: 64'b0111001011110111101001111111000010100101111101000110111111010011;
		8'd169: 64'b1010110110111011000110111011001000000011111001111100111111111010;
		8'd170: 64'b0111110011101111100000001111111111101111111111111001111110011010;
		8'd171: 64'b0110001110111011111001001010101101110101101010111101011111101011;
		8'd172: 64'b0111111100001010000100001110101101100100010110011001111100101000;
		8'd173: 64'b0011110100110101011010111011011000110111111001110010101011110110;
		8'd174: 64'b1101100111111110001111101101111111111001101101101101111011010011;
		8'd175: 64'b0101011010010000010001111100100001011000101100100111111111101010;
		8'd176: 64'b1100111101010110010110100011011101001010010110100111111010110101;
		8'd177: 64'b1100100001010111101001100100011110001100010010111011110001101001;
		8'd178: 64'b0110011101101011000111110110001011011011011010110101111111111011;
		8'd179: 64'b1011111111011110110110001010110110101010110110100100101000000111;
		8'd180: 64'b0010111011100110111111111101111100101011100101011111111101010101;
		8'd181: 64'b0010010101100111110011010101110110111101011001110110101011010000;
		8'd182: 64'b1110111101111001101011010011101100011111011110010010110110111101;
		8'd183: 64'b0011001111101111011101111100111111101111101010101111111101111010;
		8'd184: 64'b1100101111111111000110111011101011011101111011101011101111000011;
		8'd185: 64'b1101001101111001111101111111110110110111011111111111101110110101;
		8'd186: 64'b0001010101000110011111101111100000110101111001101111010111110100;
		8'd187: 64'b0001011110011000111110011011101110111111011111010011100110111011;
		8'd188: 64'b1011111010111110101010001111111110111111101001101011101110111111;
		8'd189: 64'b1111111101100010001110110110011101110001011001101101101111110110;
		8'd190: 64'b0100101111010011000101000011011101001011000111110100101111010010;
		8'd191: 64'b0101100101101100011101000111111101110011111011000111100101110110;
		8'd192: 64'b1100111101100111000011011110100111111111010100110011101111100001;
		8'd193: 64'b1110011001001011111111011011010011111111100010110111001101110111;
		8'd194: 64'b1110111110001101011101111001110111011111110011011111111011111011;
		8'd195: 64'b1111011111110111110001111111011111010111111100011101011010011111;
		8'd196: 64'b1110111010101111011111101011011100111110001001110010110111110111;
		8'd197: 64'b1111100001001101111010111011111111111100011111111011101100111110;
		8'd198: 64'b0111010001101101101011101011000101110010100011110011101010100001;
		8'd199: 64'b1010101111111011001011001110110110111101100111111100100011011110;
		8'd200: 64'b0101111101111100110101010111110111001100101111011101011101101001;
		8'd201: 64'b1010101110111110001100110010111110111011001111000011001000101011;
		8'd202: 64'b1000001110110111111101111111111111011110100001111011010110000101;
		8'd203: 64'b1011111110101111111110111110111110101001101111110001101111001010;
		8'd204: 64'b1010000110111111111001001111110011101011111101101010011100101110;
		8'd205: 64'b1111011011011000111101110001011111110110110101110100001110011101;
		8'd206: 64'b1111100010101110101011011101110100111011111011001010111011111110;
		8'd207: 64'b0111111101010111111110110111111110010101111110111111101101111111;
		8'd208: 64'b0111011010101010010010100011011111101110011110101111101001000110;
		8'd209: 64'b0110110010101111111000010010100001100000101011101010110110111100;
		8'd210: 64'b0111011111100011010111110110111111110111011001111001110101101000;
		8'd211: 64'b1111010010111110101101011111110110110000010111100111111101001100;
		8'd212: 64'b0000011111100000011111011110100011110111011000010100001011000110;
		8'd213: 64'b1011100100110011111111110111010010110011011101011011111001110100;
		8'd214: 64'b1101111111101011101111110101111110110110011011101111101101111111;
		8'd215: 64'b1110001111001100100010111011001111011101110101111000000110110001;
		8'd216: 64'b0111011001000111111001110000010100000110010010111011111101100110;
		8'd217: 64'b1111111001001010011100100010101001010011010001100111010011000011;
		8'd218: 64'b0111101111011101111110011011111010110001110101011111110111010101;
		8'd219: 64'b1010111101111101110101010111101100100101011100011100011100011101;
		8'd220: 64'b0111011011001110101101011110011101110111010101010111000110001111;
		8'd221: 64'b0001101111111001111101111101100111011111111110011101000101111111;
		8'd222: 64'b1001111000100001111111010010110100111100100100010000110110111111;
		8'd223: 64'b1111101111010111101011111100000111001001110101110100111111101001;
		8'd224: 64'b1101111011111100101011101110001011111110111111011110111001111110;
		8'd225: 64'b1010101010101011101000000010111011101111001010111111100010111110;
		8'd226: 64'b0111010101000100010110111100010101111111011101101001001111100110;
		8'd227: 64'b0010011111101001011111110011111101111101001010001011101100101111;
		8'd228: 64'b1100010010101101110101111101111111100110110111101001111100111100;
		8'd229: 64'b0101101101011000010110011101001101110011111111000001110111010110;
		8'd230: 64'b1101111111011100101011110101101000011101110110011111111011110001;
		8'd231: 64'b1001111110111001110101110100001110011011010100011001111110000001;
		8'd232: 64'b0001011110011010110101110111110100000010010111101101010011010111;
		8'd233: 64'b1111111101001010010001111010111001011111001010100111000001111110;
		8'd234: 64'b1111011011111011101011001110001111111100111110111110100100110111;
		8'd235: 64'b0111110100111000011110100101001101111100010100011111011011000100;
		8'd236: 64'b0010101111000011100110101011101010100110000011111101101100111000;
		8'd237: 64'b1010111111010111101011111000001110001011110101101101011111010111;
		8'd238: 64'b1101111011111000011100000101110111100111111111001111110011111100;
		8'd239: 64'b0111011010110011101100011111111111100001001100011000010000111111;
		8'd240: 64'b1111111111101111111101010111110111111010111011001110000111111101;
		8'd241: 64'b1111111111000111111001100101011111111010110011111110110000111100;
		8'd242: 64'b0011101110111010110001111100111110100110110010111010010111001111;
		8'd243: 64'b1111111011110101001011101011100111101100111101111101010110110001;
		8'd244: 64'b0110101111001110000000101111110100101111110011110010101010111110;
		8'd245: 64'b0010000010100111001010011111011010111101111001011111100111001100;
		8'd246: 64'b0100110101001100110011011111110001111100011110110100110111111111;
		8'd247: 64'b1100100101110101010110110011101100010011011110010010101001110101;
		8'd248: 64'b1111110001101101011111110111111011010101101111011011101111011101;
		8'd249: 64'b1110000111010110110001100010000011001010010101100101011110111111;
		8'd250: 64'b0111111100111110111111100001111111111101100111001101110100101101;
		8'd251: 64'b0101100110011111010101100101011011001110110111110111111001010110;
		8'd252: 64'b1011101001110010111110011000010111011010001100100011100110010111;
		8'd253: 64'b1001011000011101110010011101110111110001011111101001100011111110;
		8'd254: 64'b0111111111111011011110101111011110010110111110010111101101111000;
		8'd255: 64'b0101000011010101000101010111110111110001011110011101010101110101;
	endcase;
	return out;
endfunction
function Bit#(64) get_output_page6(UInt#(8) counter);
	Bit#(64) out = case(counter)
		8'd0: 64'b1111111111011011111111111101001110111110110110111011111011001000;
		8'd1: 64'b0110111010111110101010011010001011111010111100100010101111100110;
		8'd2: 64'b0011111000100010111011100111111001101011011111110110111100111111;
		8'd3: 64'b1011011011110011001101101001101010111011111111111011001111111101;
		8'd4: 64'b1101001111110011000111111110100111010011111010010111111111101000;
		8'd5: 64'b0101101011111110110110011101011110111010101110101001111111110111;
		8'd6: 64'b0101110111011101101101111110100110111100110011010111010111010101;
		8'd7: 64'b1011111111010101011111111001000111111011100110011101101111011101;
		8'd8: 64'b0101011100111011100110110110101101111111111100010101111100111011;
		8'd9: 64'b0101011110000110101110101000011111000010100011111100101010011100;
		8'd10: 64'b1111110110011100111111001111111110111111001011010011100101101100;
		8'd11: 64'b1001111101110001000111010011011000110101011101111111100110011111;
		8'd12: 64'b1010110101110111111001110111111001100111101101001111111101111010;
		8'd13: 64'b1110111011100110111100011101101000111111110010011011100110111010;
		8'd14: 64'b1101101011010110101011100111011111111110011101111110101011110101;
		8'd15: 64'b0110111100100011111101001010001111110111101101111110011111001011;
		8'd16: 64'b1010011011111111101001111111001111110111111111111111101111010001;
		8'd17: 64'b1110101111100111101001000101111111111010111001110011011001000111;
		8'd18: 64'b1010011110001001111111100110001000111011001010001110011000101010;
		8'd19: 64'b0101111010111111101111111111101111011110111110111011111110101011;
		8'd20: 64'b1011111111011101101111101111101101101111111101111111111111011111;
		8'd21: 64'b1111111111111011111111111111101111101111111110111011111111111111;
		8'd22: 64'b0110100111111010011101100110110001101101011110000011000001101001;
		8'd23: 64'b1011111010011010100011111011110111111111111010011110111110111011;
		8'd24: 64'b1111010111111111110110011011111110001101101101111111110111010111;
		8'd25: 64'b1111111111110111111110111111011110111111111101111110000101110101;
		8'd26: 64'b0001001010011111000001111111111111001111110111111000010010011111;
		8'd27: 64'b0010010111011111011010110010000100101111110011110101111111000111;
		8'd28: 64'b1100101100110010101110100101111110101011111111101000001111100110;
		8'd29: 64'b0111011111101001111111011111111111110001011111011111000111111110;
		8'd30: 64'b0101110010001011001111100100101111111010010001010001110001111001;
		8'd31: 64'b0001101110101110111110111110011101111110101001101111111111111100;
		8'd32: 64'b0101011111111100111100011111110011010011111111111001110111011000;
		8'd33: 64'b1011001101110111011001001110011100100101011101011110101101101110;
		8'd34: 64'b1011110110111110110100110110111110111010111111101111000001111111;
		8'd35: 64'b1011101111111011101111101001110110111100101111111011111110010001;
		8'd36: 64'b1101001101110011111111111111111110011111011110110111111101111111;
		8'd37: 64'b1110111111000011110111111111111111111011110010111111101111010111;
		8'd38: 64'b1101101011101111111111001111111011101111110011101111100111011110;
		8'd39: 64'b1011101111101100111111110001110100110011100010111111111100100001;
		8'd40: 64'b1110110101111110011011101111110011101101110111011100110011111100;
		8'd41: 64'b0011010101011110100111110011101010010100010111001001110000000010;
		8'd42: 64'b1100111101011011111001100101111011100111010100111110011101100111;
		8'd43: 64'b1101101111110101110111011111010110111000101101001101010101011100;
		8'd44: 64'b1111011111011101111101111011111011010111110101110011011111111110;
		8'd45: 64'b1111101111110011110011111011111111000111101110011110111111110111;
		8'd46: 64'b0100110100000100011101111111110100001101001001010100101111101100;
		8'd47: 64'b1110101101111101111011101100110011001100101101100110111011110100;
		8'd48: 64'b1111111111101111011111111101110111111011111011111110111111111111;
		8'd49: 64'b1110101110010011111011100011010111100010110100110110111100110111;
		8'd50: 64'b1000100110001111001000111100111101101111101111011011010101111111;
		8'd51: 64'b1111111010100111101111111001011010111101111011111111110011001111;
		8'd52: 64'b1111010011011110100101010111011111010111010001111100111111010111;
		8'd53: 64'b0111000100010100111101111001110000110011110110001011111011110101;
		8'd54: 64'b1111001111110111111110110101110101111011111111011111011101111011;
		8'd55: 64'b1110011011000111111001001111011010010110111101101100011111110011;
		8'd56: 64'b0110111111010101011111010111000111110101100111000111110111111011;
		8'd57: 64'b0110101101111111011101110110011101100011010111111110111101011100;
		8'd58: 64'b1110001011101111011101110100010011110111011101110110111011001101;
		8'd59: 64'b1110010000111001101111111111011111111110111110011011011111011111;
		8'd60: 64'b1101111110100101011011111111010111001111100001011110011111111101;
		8'd61: 64'b1101110100111101110111010111111111011111111101111111111111110111;
		8'd62: 64'b0111111011100110101101101001001011111010010001101111001101110111;
		8'd63: 64'b1010110011110100111101111011110001111110111110001111111111101110;
		8'd64: 64'b0100010111111111110111000101010100001101111111011101110001111011;
		8'd65: 64'b1111100111111101100110101111100110111111110111111011101110111001;
		8'd66: 64'b0111111110111010011100110111111000111010101010100111010111111111;
		8'd67: 64'b1111111100010111001111110111010101101110011101111111110110010111;
		8'd68: 64'b1011101011100110111111111111110111111111000111101100011111011111;
		8'd69: 64'b1100011101111110110101110111001011101111101101100110101100110010;
		8'd70: 64'b1001111111100100111111000111000110111101110101010101110000101011;
		8'd71: 64'b1111111110111101011110110001111011110111010111100101101110111100;
		8'd72: 64'b1110000100110111111000111001111010000101000100011100011110001110;
		8'd73: 64'b1000110111001101111111101100111110011101111011011111110011000101;
		8'd74: 64'b1111110101111001110011111101101111111111111110011111110101011111;
		8'd75: 64'b0001110011111100011111111111100001000000100111001001100011011111;
		8'd76: 64'b1110110101011110100111111011111111111101110111110011111111111001;
		8'd77: 64'b0110010100011111100010001101111100011100111111110011111111111101;
		8'd78: 64'b1010011111111111101111110111111100010101010010101111110101011011;
		8'd79: 64'b0111100010001111110011111011101101100101101011010101011010111111;
		8'd80: 64'b1111010111110101010111110111110101011100011111111101011111111101;
		8'd81: 64'b1111111010100110101011111101101011111100100011111011010110001001;
		8'd82: 64'b1100100101100010001100000000101011011101111000110111101101101010;
		8'd83: 64'b1110101101100111100111010110010101111011110001110001101111000100;
		8'd84: 64'b1011001011001110100111111110011110111110110001111011111111101111;
		8'd85: 64'b1101011100111101100111110111101100000111110001110011011111010011;
		8'd86: 64'b1111111101110111110011110111011111110111111111101111011101110101;
		8'd87: 64'b1001000011110011110110111101000111011001110110011011011110111101;
		8'd88: 64'b1000111111011111100111011101011110001110101111111000110111011101;
		8'd89: 64'b1111101110110101111100111011111110110111001100111110000101011010;
		8'd90: 64'b1111000111001111111110101101110111111100111111110111011111101111;
		8'd91: 64'b0111100000101110000111100111010100111001011001000001000010110111;
		8'd92: 64'b1110101111111010011011101111101100101111111111101110101111111011;
		8'd93: 64'b0100111110011111011110011111110111101101110111110110101111111111;
		8'd94: 64'b0111101111001101011110011111111001111111111011000100111101101010;
		8'd95: 64'b1101010111110101111100101000111111110011110101011111111001111100;
		8'd96: 64'b0010011111101011111110111110111100111101111111110011111111101101;
		8'd97: 64'b1011111110101010111111111011100010110111101010101111111011101101;
		8'd98: 64'b1110001100111011101011111001101101110011001100100111011000110111;
		8'd99: 64'b0111110111110111011001101111000111010101101101101110010111100100;
		8'd100: 64'b1101111100011001111111011110101111011101101110011101001111111100;
		8'd101: 64'b0011100100100000010001001111011101011011101001110101011110010110;
		8'd102: 64'b0101110011011111111111111111111111111110111111111101111001010111;
		8'd103: 64'b0111011101010011001010111010001011110011011110100110001111010110;
		8'd104: 64'b1110111110011011111100011000111111010011011010111111110111111011;
		8'd105: 64'b0110011011000111011101110010111100101111001111110111110100111011;
		8'd106: 64'b1010111110111011011111101011111110101111011100110010111111111001;
		8'd107: 64'b1011110110111001010011110111100010010011001110010010111001100001;
		8'd108: 64'b1111111100101111011111110111011111011111010011111111111101111111;
		8'd109: 64'b0101111010100110000111111111111011001010111001110110111100110111;
		8'd110: 64'b0110011011111111011001011010110101101101001111010111011011110101;
		8'd111: 64'b0111001111111111111110010111011111111111101011101110111101110110;
		8'd112: 64'b1101100001011111111111100011010011111100110101111111111011110101;
		8'd113: 64'b1011011000001111111111001110100110110011000111001011111110101000;
		8'd114: 64'b1101001000011011001100110010000110011101010111011111011001111011;
		8'd115: 64'b0111101111100101011111111110111101110111111001000010111111111111;
		8'd116: 64'b1011111110101111101111010011100111011101000001011011111100111001;
		8'd117: 64'b0111101100101011101010111110111101001110111001111010111011110111;
		8'd118: 64'b1110111111010111001011001111011001010111110011100010111001000100;
		8'd119: 64'b0111011101111111111100111000001111010111011111001101010101000011;
		8'd120: 64'b0111001111111111110101010111001111100111011111110010011001111111;
		8'd121: 64'b0101101111111111001110100001001111011110011111000001100100111101;
		8'd122: 64'b1011010111011101110110101001101010010011111110111001101101011011;
		8'd123: 64'b0011001001010010101100101000000101101111010101100110101111001010;
		8'd124: 64'b1100101101001100111001111011010011001100011011111110101011101111;
		8'd125: 64'b1011010010111011101010001100110010100100110111101011010110111011;
		8'd126: 64'b0111111011001011001111110001101010110111011001111011011010011011;
		8'd127: 64'b0111111110110111100110111010110100100110111101010101000101100111;
		8'd128: 64'b1100110001111111111111111111110011101111111011111110111111111111;
		8'd129: 64'b1111101111001111111011101110111111111010111011111110011101011110;
		8'd130: 64'b1101000111000111011011111000110111111101100011110101111111100111;
		8'd131: 64'b1100001010110010011001101101100011010111111011111110111110010011;
		8'd132: 64'b1111000110111111110011100110011111001111011111111000111001100110;
		8'd133: 64'b0100001011000111111111001111110101011011110111110111111111011111;
		8'd134: 64'b1011011011111111111101011101110111110011011011110101111111011111;
		8'd135: 64'b1100111010110101111100111111100110111010101011001111110111010010;
		8'd136: 64'b0011111110111111101111111011111111101111000111111011110111111111;
		8'd137: 64'b1001100110111111010010111111111101011001101110101100110100111011;
		8'd138: 64'b0011101110110110001011001101110000111001101011100010100100111110;
		8'd139: 64'b1001111000001111110111101000110110011101011011011110111101111101;
		8'd140: 64'b0111101011101110100101100101101100101010010100101101111011110111;
		8'd141: 64'b1001010011000001110100111110111011110110110001010000111011001100;
		8'd142: 64'b1101111010101110111111111010101010011111101111001011100010101010;
		8'd143: 64'b1111101000111010101101000011001111110011010010100010001001010111;
		8'd144: 64'b0100100110001001011001110110100110100111111110010101101100111110;
		8'd145: 64'b0101101001111011111111111011101100110011001110101111101101110011;
		8'd146: 64'b1011101111111111111101101101101111000001100110111011011001001111;
		8'd147: 64'b0111111101101111010110101111111111110111111111110100111110111111;
		8'd148: 64'b1100001101101010010000111011000001011001011010000100010101011111;
		8'd149: 64'b1111111111101111010111101110011111100111111011111101011011001111;
		8'd150: 64'b1010111010011110101111111110111010111111111010001010111011111111;
		8'd151: 64'b1010111010011111101011101000110110101010100011111110101110001011;
		8'd152: 64'b1111010101111011011011111111101000111101001111111111101101111010;
		8'd153: 64'b1011011011001000011101111010011011110011111111100111111101111010;
		8'd154: 64'b1101111111101110100111111111111110011111111111111001111110111101;
		8'd155: 64'b1101111110110111111101111011110111111011101101010011011110110101;
		8'd156: 64'b1010111010011110111110111111110100101110110110001000110111001111;
		8'd157: 64'b0010101110001011110011101010011110010000001001111110110110001100;
		8'd158: 64'b0111111000011111011001110111111110100110001111101010011000101111;
		8'd159: 64'b1111011110110111110101101001011110110111111101111011011010101011;
		8'd160: 64'b0111101111111111111010111111111101111101111101101111101011111111;
		8'd161: 64'b0111100110111001111101100010110011011111101011111001101100011100;
		8'd162: 64'b1111101111111111011101011110011101111111111101111110101011100111;
		8'd163: 64'b1001000101111101101110111000101111101001101110011110100101001101;
		8'd164: 64'b1111101110101111101110111110110010111111111011100010100111111100;
		8'd165: 64'b0001010000110110011101110010111100011010101011101001001110111111;
		8'd166: 64'b1011001111010111001101110111001110100101111111110011111101010111;
		8'd167: 64'b1101101111100011111101101111011111010111111100011111011011100111;
		8'd168: 64'b0111011011110111101001111111000011100101111101000110111111010011;
		8'd169: 64'b1010111110111011000110111011111000000111111001111100111111111010;
		8'd170: 64'b0111110011101111100000001111111111111111111111111001111110011110;
		8'd171: 64'b0110001110111011111001001010101101110101101010111101011111101011;
		8'd172: 64'b0111111100001010000111001110101101110100010110011001111100101000;
		8'd173: 64'b0011110100110111011011111011011100110111111001110010101011111110;
		8'd174: 64'b1101100111111110001111101101111111111011101101101101111011010011;
		8'd175: 64'b0101011010110000010011111101100001011000101100100111111111101010;
		8'd176: 64'b1100111101010110010111100111011101001010010110100111111010110101;
		8'd177: 64'b1100100001010111101011100110111110001100010010111011110001101001;
		8'd178: 64'b0110011101101011000111110110001011011011011110110101111111111011;
		8'd179: 64'b1011111111011110110110001010110111101110110110110100101000000111;
		8'd180: 64'b0110111011100111111111111111111100101011110101011111111101010101;
		8'd181: 64'b0110010101100111111011010101110110111101011011111110101011010010;
		8'd182: 64'b1110111101111001101011010011101110011111011110010011110110111101;
		8'd183: 64'b0011001111101111011101111111111111101111101011101111111101111010;
		8'd184: 64'b1100101111111111101110111011101011011101111011111011101111000011;
		8'd185: 64'b1101001101111001111101111111110110110111011111111111101110110101;
		8'd186: 64'b0001010101000110011111101111101000110101111001101111010111110100;
		8'd187: 64'b0011011110011000111110011011101110111111011111010011100110111011;
		8'd188: 64'b1111111010111110101010101111111110111111101001101011111110111111;
		8'd189: 64'b1111111101100010011110110110011101110001011101101101101111110110;
		8'd190: 64'b0100101111010011000101000011111101001011000111110101101111010010;
		8'd191: 64'b0101100101101100011101000111111101110011111111000111110101110111;
		8'd192: 64'b1100111101100111000011011110100111111111010100110011101111100001;
		8'd193: 64'b1110011001001011111111011011010011111111100010110111001101110111;
		8'd194: 64'b1111111110001101011101111001110111011111110111111111111111111011;
		8'd195: 64'b1111011111110111110001111111011111010111111100011101011010011111;
		8'd196: 64'b1110111010101111011111111111011110111110111101110010110111110111;
		8'd197: 64'b1111100001001101111011111011111111111100011111111011101100111110;
		8'd198: 64'b1111010001101101101011111011000101110010101011110011101010100001;
		8'd199: 64'b1010101111111011101011001110110111111101100111111100100011111110;
		8'd200: 64'b0101111101111100110101010111110111001100101111011101011101101001;
		8'd201: 64'b1010101110111110101110110011111110111011001111000011001000101011;
		8'd202: 64'b1000001110110111111101111111111111011110100001111011010110000101;
		8'd203: 64'b1011111110101111111110111110111110101001101111110001101111001010;
		8'd204: 64'b1110000110111111111001001111111011101011111101101010011110111110;
		8'd205: 64'b1111011011011000111101110001011111110110110101110101011110011101;
		8'd206: 64'b1111101010101110101011011101110100111111111011001011111011111110;
		8'd207: 64'b0111111101010111111110110111111111110101111110111111101101111111;
		8'd208: 64'b0111011010101010010010100011011111101110111110101111101001000110;
		8'd209: 64'b0110110010101111111000010010100001100000101011101010110110111100;
		8'd210: 64'b1111011111101011011111110110111111111111011101111001110101101000;
		8'd211: 64'b1111010010111110101101011111110110110010010111100111111101001101;
		8'd212: 64'b0000011111110010011111111110100011110111011000011100001011010110;
		8'd213: 64'b1011100101110011111111111111010010111011011101011011111101110100;
		8'd214: 64'b1101111111101011101111110101111110110111111011111111111101111111;
		8'd215: 64'b1111001111011100100010111011001111011101110101111000000110110101;
		8'd216: 64'b0111011001100111111001110010010100000110010010111011111111100110;
		8'd217: 64'b1111111001001010011100100011101011010111110011100111011011000111;
		8'd218: 64'b0111101111011111111110011011111011110001110101011111110111010101;
		8'd219: 64'b1010111101111101110101010111101100100101011100011100011100011101;
		8'd220: 64'b0111011011001110101101011110111101110111010101010111000110101111;
		8'd221: 64'b0001101111111001111101111101100111011111111110011101000111111111;
		8'd222: 64'b1001111000100001111111010010110100111100100100010001110111111111;
		8'd223: 64'b1111101111010111111011111101000111111001110101110100111111101001;
		8'd224: 64'b1101111011111111111011101110001111111110111111011110111001111110;
		8'd225: 64'b1010101010101011101000000010111011101111001010111111100010111110;
		8'd226: 64'b0111010101000110010110111100010101111111011101111001001111101110;
		8'd227: 64'b0010011111101001011111110111111101111101001010011011111100101111;
		8'd228: 64'b1100010010101101110101111101111111100110110111101001111100111100;
		8'd229: 64'b0101101101011100010110011101001101110011111111101001110111010111;
		8'd230: 64'b1101111111011100101011110101101000011101110110011111111011110001;
		8'd231: 64'b1001111110111001110111110110001110011011010100011001111110000001;
		8'd232: 64'b0101011110011110110101111111110100000010110111101101010111010111;
		8'd233: 64'b1111111101001010010001111010111001011111011010100111000001111110;
		8'd234: 64'b1111011011111011101011001110001111111100111110111110100100110111;
		8'd235: 64'b0111110100111000011110100101001101111100010100011111011111000100;
		8'd236: 64'b0010101111000111100110101011101010100110000011111101101110111010;
		8'd237: 64'b1010111111110111101011111000101110101011110101101101011111010111;
		8'd238: 64'b1101111011111000011100000101110111110111111111001111110011111100;
		8'd239: 64'b0111011010110111101100011111111111100001001100111000010000111111;
		8'd240: 64'b1111111111101111111101011111111111111010111011011111000111111101;
		8'd241: 64'b1111111111010111111001100101011111111010110011111110110001111100;
		8'd242: 64'b1011101110111010110001111100111110100110110010111010110111001111;
		8'd243: 64'b1111111011110101001011101011100111101100111101111101010110110001;
		8'd244: 64'b0110111111001110000000101111110100111111110011110010101011111110;
		8'd245: 64'b0010000010100111001010011111011010111101111001011111100111001100;
		8'd246: 64'b0110110101001100110011011111110001111100011110110100110111111111;
		8'd247: 64'b1100100101110101010110110011101100010011011110010010101001110101;
		8'd248: 64'b1111110011101101011111110111111011011101111111011011101111011101;
		8'd249: 64'b1110000111010110110001100011000011011010010101100101011110111111;
		8'd250: 64'b0111111100111110111111100011111111111101100111111101110100111101;
		8'd251: 64'b0101100110011111010101100101011011001110110111110111111001010110;
		8'd252: 64'b1011101001110011111110011001010111011010001100100011100110010111;
		8'd253: 64'b1101011000011101110010011101110111110001011111101001100011111110;
		8'd254: 64'b0111111111111011011110101111011111010110111110010111101101111000;
		8'd255: 64'b0101010111010101010101010111110111110001011110011101010101110101;
	endcase;
	return out;
endfunction
